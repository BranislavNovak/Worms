
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity ram is
	generic
	(
		DATA_WIDTH : natural := 32;		    -- 4 byte one line of memory
		ADDR_WIDTH : natural := 13			    -- 24576 bytes size of memory
	);

	port(
		i_clk    : in  std_logic;
		i_r_addr : in  std_logic_vector(ADDR_WIDTH-1 downto 0);
		i_data   : in  std_logic_vector(DATA_WIDTH-1 downto 0);
		i_we     : in  std_logic;
		i_w_addr : in  std_logic_vector(ADDR_WIDTH-1 downto 0);
		o_data   : out std_logic_vector(DATA_WIDTH-1 downto 0)
	);
end entity ram;

architecture arch of ram is

	type ram_t is array (0 to 2**ADDR_WIDTH-1) of std_logic_vector(DATA_WIDTH-1 downto 0);


-- GENERATED BY BC_MEM_PACKER

-- DATE: Thu May 18 16:01:02 2017

	signal mem : ram_t := (

--			***** COLOR PALLETE *****


		0 =>	x"01010101", -- R: 0 G: 0 B: 0
		1 =>	x"00FFFFFF", -- R: 255 G: 255 B: 255
		2 =>	x"00F0FBFF", -- R: 255 G: 251 B: 240
		3 =>	x"00C0C0C0", -- R: 192 G: 192 B: 192
		4 =>	x"00C0DCC0", -- R: 192 G: 220 B: 192
		5 =>	x"00404040", -- R: 64 G: 64 B: 64
		6 =>	x"00808080", -- R: 128 G: 128 B: 128
		7 =>	x"0080A0A0", -- R: 160 G: 160 B: 128
		8 =>	x"00406080", -- R: 128 G: 96 B: 64
		9 =>	x"008080A0", -- R: 160 G: 128 B: 128
		10 =>	x"008080C0", -- R: 192 G: 128 B: 128
		11 =>	x"004060A0", -- R: 160 G: 96 B: 64
		12 =>	x"0080A0E0", -- R: 224 G: 160 B: 128
		13 =>	x"0080A0C0", -- R: 192 G: 160 B: 128
		14 =>	x"008080E0", -- R: 224 G: 128 B: 128
		15 =>	x"008060C0", -- R: 192 G: 96 B: 128
		16 =>	x"008060E0", -- R: 224 G: 96 B: 128
		17 =>	x"0080C0E0", -- R: 224 G: 192 B: 128
		18 =>	x"00A4A0A0", -- R: 160 G: 160 B: 164
		19 =>	x"00808060", -- R: 96 G: 128 B: 128
		20 =>	x"00806060", -- R: 96 G: 96 B: 128
		21 =>	x"0080A080", -- R: 128 G: 160 B: 128
		22 =>	x"00C0A080", -- R: 128 G: 160 B: 192
		23 =>	x"00C0A060", -- R: 96 G: 160 B: 192
		24 =>	x"00806040", -- R: 64 G: 96 B: 128
		25 =>	x"00806020", -- R: 32 G: 96 B: 128
		26 =>	x"00406060", -- R: 96 G: 96 B: 64
		27 =>	x"00004080", -- R: 128 G: 64 B: 0
		28 =>	x"00404060", -- R: 96 G: 64 B: 64
		29 =>	x"00006080", -- R: 128 G: 96 B: 0
		30 =>	x"00004060", -- R: 96 G: 64 B: 0
		31 =>	x"00002040", -- R: 64 G: 32 B: 0
		32 =>	x"00404080", -- R: 128 G: 64 B: 64
		33 =>	x"004060C0", -- R: 192 G: 96 B: 64
		34 =>	x"00C0A000", -- R: 0 G: 160 B: 192
		35 =>	x"008060A0", -- R: 160 G: 96 B: 128
		36 =>	x"00002060", -- R: 96 G: 32 B: 0
		37 =>	x"004080A0", -- R: 160 G: 128 B: 64
		38 =>	x"00402060", -- R: 96 G: 32 B: 64
		39 =>	x"004080C0", -- R: 192 G: 128 B: 64
		40 =>	x"00000000", -- Unused
		41 =>	x"00000000", -- Unused
		42 =>	x"00000000", -- Unused
		43 =>	x"00000000", -- Unused
		44 =>	x"00000000", -- Unused
		45 =>	x"00000000", -- Unused
		46 =>	x"00000000", -- Unused
		47 =>	x"00000000", -- Unused
		48 =>	x"00000000", -- Unused
		49 =>	x"00000000", -- Unused
		50 =>	x"00000000", -- Unused
		51 =>	x"00000000", -- Unused
		52 =>	x"00000000", -- Unused
		53 =>	x"00000000", -- Unused
		54 =>	x"00000000", -- Unused
		55 =>	x"00000000", -- Unused
		56 =>	x"00000000", -- Unused
		57 =>	x"00000000", -- Unused
		58 =>	x"00000000", -- Unused
		59 =>	x"00000000", -- Unused
		60 =>	x"00000000", -- Unused
		61 =>	x"00000000", -- Unused
		62 =>	x"00000000", -- Unused
		63 =>	x"00000000", -- Unused
		64 =>	x"00000000", -- Unused
		65 =>	x"00000000", -- Unused
		66 =>	x"00000000", -- Unused
		67 =>	x"00000000", -- Unused
		68 =>	x"00000000", -- Unused
		69 =>	x"00000000", -- Unused
		70 =>	x"00000000", -- Unused
		71 =>	x"00000000", -- Unused
		72 =>	x"00000000", -- Unused
		73 =>	x"00000000", -- Unused
		74 =>	x"00000000", -- Unused
		75 =>	x"00000000", -- Unused
		76 =>	x"00000000", -- Unused
		77 =>	x"00000000", -- Unused
		78 =>	x"00000000", -- Unused
		79 =>	x"00000000", -- Unused
		80 =>	x"00000000", -- Unused
		81 =>	x"00000000", -- Unused
		82 =>	x"00000000", -- Unused
		83 =>	x"00000000", -- Unused
		84 =>	x"00000000", -- Unused
		85 =>	x"00000000", -- Unused
		86 =>	x"00000000", -- Unused
		87 =>	x"00000000", -- Unused
		88 =>	x"00000000", -- Unused
		89 =>	x"00000000", -- Unused
		90 =>	x"00000000", -- Unused
		91 =>	x"00000000", -- Unused
		92 =>	x"00000000", -- Unused
		93 =>	x"00000000", -- Unused
		94 =>	x"00000000", -- Unused
		95 =>	x"00000000", -- Unused
		96 =>	x"00000000", -- Unused
		97 =>	x"00000000", -- Unused
		98 =>	x"00000000", -- Unused
		99 =>	x"00000000", -- Unused
		100 =>	x"00000000", -- Unused
		101 =>	x"00000000", -- Unused
		102 =>	x"00000000", -- Unused
		103 =>	x"00000000", -- Unused
		104 =>	x"00000000", -- Unused
		105 =>	x"00000000", -- Unused
		106 =>	x"00000000", -- Unused
		107 =>	x"00000000", -- Unused
		108 =>	x"00000000", -- Unused
		109 =>	x"00000000", -- Unused
		110 =>	x"00000000", -- Unused
		111 =>	x"00000000", -- Unused
		112 =>	x"00000000", -- Unused
		113 =>	x"00000000", -- Unused
		114 =>	x"00000000", -- Unused
		115 =>	x"00000000", -- Unused
		116 =>	x"00000000", -- Unused
		117 =>	x"00000000", -- Unused
		118 =>	x"00000000", -- Unused
		119 =>	x"00000000", -- Unused
		120 =>	x"00000000", -- Unused
		121 =>	x"00000000", -- Unused
		122 =>	x"00000000", -- Unused
		123 =>	x"00000000", -- Unused
		124 =>	x"00000000", -- Unused
		125 =>	x"00000000", -- Unused
		126 =>	x"00000000", -- Unused
		127 =>	x"00000000", -- Unused
		128 =>	x"00000000", -- Unused
		129 =>	x"00000000", -- Unused
		130 =>	x"00000000", -- Unused
		131 =>	x"00000000", -- Unused
		132 =>	x"00000000", -- Unused
		133 =>	x"00000000", -- Unused
		134 =>	x"00000000", -- Unused
		135 =>	x"00000000", -- Unused
		136 =>	x"00000000", -- Unused
		137 =>	x"00000000", -- Unused
		138 =>	x"00000000", -- Unused
		139 =>	x"00000000", -- Unused
		140 =>	x"00000000", -- Unused
		141 =>	x"00000000", -- Unused
		142 =>	x"00000000", -- Unused
		143 =>	x"00000000", -- Unused
		144 =>	x"00000000", -- Unused
		145 =>	x"00000000", -- Unused
		146 =>	x"00000000", -- Unused
		147 =>	x"00000000", -- Unused
		148 =>	x"00000000", -- Unused
		149 =>	x"00000000", -- Unused
		150 =>	x"00000000", -- Unused
		151 =>	x"00000000", -- Unused
		152 =>	x"00000000", -- Unused
		153 =>	x"00000000", -- Unused
		154 =>	x"00000000", -- Unused
		155 =>	x"00000000", -- Unused
		156 =>	x"00000000", -- Unused
		157 =>	x"00000000", -- Unused
		158 =>	x"00000000", -- Unused
		159 =>	x"00000000", -- Unused
		160 =>	x"00000000", -- Unused
		161 =>	x"00000000", -- Unused
		162 =>	x"00000000", -- Unused
		163 =>	x"00000000", -- Unused
		164 =>	x"00000000", -- Unused
		165 =>	x"00000000", -- Unused
		166 =>	x"00000000", -- Unused
		167 =>	x"00000000", -- Unused
		168 =>	x"00000000", -- Unused
		169 =>	x"00000000", -- Unused
		170 =>	x"00000000", -- Unused
		171 =>	x"00000000", -- Unused
		172 =>	x"00000000", -- Unused
		173 =>	x"00000000", -- Unused
		174 =>	x"00000000", -- Unused
		175 =>	x"00000000", -- Unused
		176 =>	x"00000000", -- Unused
		177 =>	x"00000000", -- Unused
		178 =>	x"00000000", -- Unused
		179 =>	x"00000000", -- Unused
		180 =>	x"00000000", -- Unused
		181 =>	x"00000000", -- Unused
		182 =>	x"00000000", -- Unused
		183 =>	x"00000000", -- Unused
		184 =>	x"00000000", -- Unused
		185 =>	x"00000000", -- Unused
		186 =>	x"00000000", -- Unused
		187 =>	x"00000000", -- Unused
		188 =>	x"00000000", -- Unused
		189 =>	x"00000000", -- Unused
		190 =>	x"00000000", -- Unused
		191 =>	x"00000000", -- Unused
		192 =>	x"00000000", -- Unused
		193 =>	x"00000000", -- Unused
		194 =>	x"00000000", -- Unused
		195 =>	x"00000000", -- Unused
		196 =>	x"00000000", -- Unused
		197 =>	x"00000000", -- Unused
		198 =>	x"00000000", -- Unused
		199 =>	x"00000000", -- Unused
		200 =>	x"00000000", -- Unused
		201 =>	x"00000000", -- Unused
		202 =>	x"00000000", -- Unused
		203 =>	x"00000000", -- Unused
		204 =>	x"00000000", -- Unused
		205 =>	x"00000000", -- Unused
		206 =>	x"00000000", -- Unused
		207 =>	x"00000000", -- Unused
		208 =>	x"00000000", -- Unused
		209 =>	x"00000000", -- Unused
		210 =>	x"00000000", -- Unused
		211 =>	x"00000000", -- Unused
		212 =>	x"00000000", -- Unused
		213 =>	x"00000000", -- Unused
		214 =>	x"00000000", -- Unused
		215 =>	x"00000000", -- Unused
		216 =>	x"00000000", -- Unused
		217 =>	x"00000000", -- Unused
		218 =>	x"00000000", -- Unused
		219 =>	x"00000000", -- Unused
		220 =>	x"00000000", -- Unused
		221 =>	x"00000000", -- Unused
		222 =>	x"00000000", -- Unused
		223 =>	x"00000000", -- Unused
		224 =>	x"00000000", -- Unused
		225 =>	x"00000000", -- Unused
		226 =>	x"00000000", -- Unused
		227 =>	x"00000000", -- Unused
		228 =>	x"00000000", -- Unused
		229 =>	x"00000000", -- Unused
		230 =>	x"00000000", -- Unused
		231 =>	x"00000000", -- Unused
		232 =>	x"00000000", -- Unused
		233 =>	x"00000000", -- Unused
		234 =>	x"00000000", -- Unused
		235 =>	x"00000000", -- Unused
		236 =>	x"00000000", -- Unused
		237 =>	x"00000000", -- Unused
		238 =>	x"00000000", -- Unused
		239 =>	x"00000000", -- Unused
		240 =>	x"00000000", -- Unused
		241 =>	x"00000000", -- Unused
		242 =>	x"00000000", -- Unused
		243 =>	x"00000000", -- Unused
		244 =>	x"00000000", -- Unused
		245 =>	x"00000000", -- Unused
		246 =>	x"00000000", -- Unused
		247 =>	x"00000000", -- Unused
		248 =>	x"00000000", -- Unused
		249 =>	x"00000000", -- Unused
		250 =>	x"00000000", -- Unused
		251 =>	x"00000000", -- Unused
		252 =>	x"00000000", -- Unused
		253 =>	x"00000000", -- Unused
		254 =>	x"00000000", -- Unused

--			***** 16x16 IMAGES *****




		255 =>	x"01010101", -- IMG_16x18_crvcina_desno
		256 =>	x"01010101",
		257 =>	x"02030101",
		258 =>	x"01010101",
		259 =>	x"01010101",
		260 =>	x"01020401",
		261 =>	x"05050101",
		262 =>	x"01010101",
		263 =>	x"01010101",
		264 =>	x"01060007",
		265 =>	x"08090101",
		266 =>	x"01010101",
		267 =>	x"01010101",
		268 =>	x"030A0B0C",
		269 =>	x"0C0D0201",
		270 =>	x"01010101",
		271 =>	x"0101010D",
		272 =>	x"0E0C0C0C",
		273 =>	x"0C0C0301",
		274 =>	x"01010101",
		275 =>	x"0101010F",
		276 =>	x"0E0E0C0C",
		277 =>	x"0E0C0301",
		278 =>	x"01010101",
		279 =>	x"0101010A",
		280 =>	x"100E0303",
		281 =>	x"0C030301",
		282 =>	x"04060201",
		283 =>	x"01010103",
		284 =>	x"0F0E0C11",
		285 =>	x"0C0C1204",
		286 =>	x"06131415",
		287 =>	x"01010101",
		288 =>	x"0D0F0912",
		289 =>	x"12121216",
		290 =>	x"17131806",
		291 =>	x"01020303",
		292 =>	x"03061913",
		293 =>	x"131A1B1C",
		294 =>	x"13131201",
		295 =>	x"01081B1D",
		296 =>	x"1B131616",
		297 =>	x"181E1B08",
		298 =>	x"1A120201",
		299 =>	x"02081B1E",
		300 =>	x"1F200A09",
		301 =>	x"1C210F0A",
		302 =>	x"03010101",
		303 =>	x"021A1F1F",
		304 =>	x"2010100E",
		305 =>	x"0C0E0A03",
		306 =>	x"01010101",
		307 =>	x"121A1F08",
		308 =>	x"0F0F0B0A",
		309 =>	x"0C0D0D02",
		310 =>	x"01010101",
		311 =>	x"01020402",
		312 =>	x"02040402",
		313 =>	x"02020101",
		314 =>	x"01010101",
		315 =>	x"01010101",
		316 =>	x"01010101",
		317 =>	x"01010101",
		318 =>	x"01010101",
		319 =>	x"01010101", -- IMG_16x18_crvcina_levo
		320 =>	x"01010302",
		321 =>	x"01010101",
		322 =>	x"01010101",
		323 =>	x"01010101",
		324 =>	x"01010505",
		325 =>	x"01040201",
		326 =>	x"01010101",
		327 =>	x"01010101",
		328 =>	x"01010908",
		329 =>	x"07000601",
		330 =>	x"01010101",
		331 =>	x"01010101",
		332 =>	x"01020D0C",
		333 =>	x"0C0B0A03",
		334 =>	x"01010101",
		335 =>	x"01010101",
		336 =>	x"01030C0C",
		337 =>	x"0C0C0C0E",
		338 =>	x"0D010101",
		339 =>	x"01010101",
		340 =>	x"01030C0E",
		341 =>	x"0C0C0E0E",
		342 =>	x"0F010101",
		343 =>	x"01020604",
		344 =>	x"0103030C",
		345 =>	x"03030E10",
		346 =>	x"0A010101",
		347 =>	x"15141306",
		348 =>	x"04120C0C",
		349 =>	x"110C0E0F",
		350 =>	x"03010101",
		351 =>	x"06181317",
		352 =>	x"16121212",
		353 =>	x"12090F0D",
		354 =>	x"01010101",
		355 =>	x"01121313",
		356 =>	x"1C1B1A13",
		357 =>	x"13190603",
		358 =>	x"03030201",
		359 =>	x"0102121A",
		360 =>	x"081B1E18",
		361 =>	x"1616131B",
		362 =>	x"1D1B0801",
		363 =>	x"01010103",
		364 =>	x"0A0F211C",
		365 =>	x"090A201F",
		366 =>	x"1E1B0802",
		367 =>	x"01010101",
		368 =>	x"030A0E0C",
		369 =>	x"0E101020",
		370 =>	x"1F1F1A02",
		371 =>	x"01010101",
		372 =>	x"020D0D0C",
		373 =>	x"0A0B0F0F",
		374 =>	x"081F1A12",
		375 =>	x"01010101",
		376 =>	x"01010202",
		377 =>	x"02040402",
		378 =>	x"02040201",
		379 =>	x"01010101",
		380 =>	x"01010101",
		381 =>	x"01010101",
		382 =>	x"01010101",
		383 =>	x"22222222", -- IMG_16x18_nebo_svetlo
		384 =>	x"22222222",
		385 =>	x"22222222",
		386 =>	x"22222222",
		387 =>	x"22222222",
		388 =>	x"22222222",
		389 =>	x"22222222",
		390 =>	x"22222222",
		391 =>	x"22222222",
		392 =>	x"22222222",
		393 =>	x"22222222",
		394 =>	x"22222222",
		395 =>	x"22222222",
		396 =>	x"22222222",
		397 =>	x"22222222",
		398 =>	x"22222222",
		399 =>	x"22222222",
		400 =>	x"22222222",
		401 =>	x"22222222",
		402 =>	x"22222222",
		403 =>	x"22222222",
		404 =>	x"22222222",
		405 =>	x"22222222",
		406 =>	x"22222222",
		407 =>	x"22222222",
		408 =>	x"22222222",
		409 =>	x"22222222",
		410 =>	x"22222222",
		411 =>	x"22222222",
		412 =>	x"22222222",
		413 =>	x"22222222",
		414 =>	x"22222222",
		415 =>	x"22222222",
		416 =>	x"22222222",
		417 =>	x"22222222",
		418 =>	x"22222222",
		419 =>	x"22222222",
		420 =>	x"22222222",
		421 =>	x"22222222",
		422 =>	x"22222222",
		423 =>	x"22222222",
		424 =>	x"22222222",
		425 =>	x"22222222",
		426 =>	x"22222222",
		427 =>	x"22222222",
		428 =>	x"22222222",
		429 =>	x"22222222",
		430 =>	x"22222222",
		431 =>	x"22222222",
		432 =>	x"22222222",
		433 =>	x"22222222",
		434 =>	x"22222222",
		435 =>	x"22222222",
		436 =>	x"22222222",
		437 =>	x"22222222",
		438 =>	x"22222222",
		439 =>	x"22222222",
		440 =>	x"22222222",
		441 =>	x"22222222",
		442 =>	x"22222222",
		443 =>	x"22222222",
		444 =>	x"22222222",
		445 =>	x"22222222",
		446 =>	x"22222222",
		447 =>	x"01010101", -- IMG_16x18_oblak
		448 =>	x"01010101",
		449 =>	x"01010101",
		450 =>	x"01010101",
		451 =>	x"01010101",
		452 =>	x"01010101",
		453 =>	x"01010101",
		454 =>	x"01010101",
		455 =>	x"01010101",
		456 =>	x"01010101",
		457 =>	x"01010101",
		458 =>	x"01010101",
		459 =>	x"01010101",
		460 =>	x"01010101",
		461 =>	x"01010101",
		462 =>	x"01010101",
		463 =>	x"01010101",
		464 =>	x"01010101",
		465 =>	x"01010101",
		466 =>	x"01010101",
		467 =>	x"01010101",
		468 =>	x"01010101",
		469 =>	x"01010101",
		470 =>	x"01010101",
		471 =>	x"01010101",
		472 =>	x"01010101",
		473 =>	x"01010101",
		474 =>	x"01010101",
		475 =>	x"01010101",
		476 =>	x"01010101",
		477 =>	x"01010101",
		478 =>	x"01010101",
		479 =>	x"01010101",
		480 =>	x"01010101",
		481 =>	x"01010101",
		482 =>	x"01010101",
		483 =>	x"01010101",
		484 =>	x"01010101",
		485 =>	x"01010101",
		486 =>	x"01010101",
		487 =>	x"01010101",
		488 =>	x"01010101",
		489 =>	x"01010101",
		490 =>	x"01010101",
		491 =>	x"01010101",
		492 =>	x"01010101",
		493 =>	x"01010101",
		494 =>	x"01010101",
		495 =>	x"01010101",
		496 =>	x"01010101",
		497 =>	x"01010101",
		498 =>	x"01010101",
		499 =>	x"01010101",
		500 =>	x"01010101",
		501 =>	x"01010101",
		502 =>	x"01010101",
		503 =>	x"01010101",
		504 =>	x"01010101",
		505 =>	x"01010101",
		506 =>	x"01010101",
		507 =>	x"01010101",
		508 =>	x"01010101",
		509 =>	x"01010101",
		510 =>	x"01010101",
		511 =>	x"0B0B0808", -- IMG_16x18_tobla1
		512 =>	x"200B2008",
		513 =>	x"0B0B2020",
		514 =>	x"20200B0B",
		515 =>	x"2020200B",
		516 =>	x"08202320",
		517 =>	x"200B0B0B",
		518 =>	x"0B202020",
		519 =>	x"200B2308",
		520 =>	x"0B0B200B",
		521 =>	x"0B202020",
		522 =>	x"20200B20",
		523 =>	x"080B080B",
		524 =>	x"0B0B2008",
		525 =>	x"080B0B0B",
		526 =>	x"2020200B",
		527 =>	x"0B0B0808",
		528 =>	x"0B23080B",
		529 =>	x"200B2020",
		530 =>	x"0B0B2024",
		531 =>	x"0B090820",
		532 =>	x"090B080B",
		533 =>	x"0B08080B",
		534 =>	x"0B0B2308",
		535 =>	x"0B202308",
		536 =>	x"0B0B0823",
		537 =>	x"0B0B0B0B",
		538 =>	x"0908080B",
		539 =>	x"0B230B0B",
		540 =>	x"0B0B0B0A",
		541 =>	x"0B0B0B0B",
		542 =>	x"0B0B0B20",
		543 =>	x"0B230820",
		544 =>	x"0B0A090B",
		545 =>	x"080A0B0A",
		546 =>	x"20080B0B",
		547 =>	x"08200B0B",
		548 =>	x"230B0A09",
		549 =>	x"0A090B0B",
		550 =>	x"0B08230B",
		551 =>	x"0B200B0B",
		552 =>	x"0B0B0B0B",
		553 =>	x"0808200B",
		554 =>	x"200B0B0B",
		555 =>	x"0B230B0B",
		556 =>	x"08200B0B",
		557 =>	x"0B250B0B",
		558 =>	x"0B0A2020",
		559 =>	x"0A200B0B",
		560 =>	x"200A0B0B",
		561 =>	x"200B0B20",
		562 =>	x"0B0A2008",
		563 =>	x"200B0B0A",
		564 =>	x"200B080B",
		565 =>	x"0B0B090B",
		566 =>	x"0B0A0B0B",
		567 =>	x"200B0A0B",
		568 =>	x"230B200B",
		569 =>	x"0B240B0B",
		570 =>	x"0B0B0B26",
		571 =>	x"0B0A2320",
		572 =>	x"0B0A0B0B",
		573 =>	x"0A0B0A0B",
		574 =>	x"0B0B0808",
		575 =>	x"27272727", -- IMG_16x18_tobla2
		576 =>	x"27272727",
		577 =>	x"27272727",
		578 =>	x"27272727",
		579 =>	x"27272727",
		580 =>	x"27272727",
		581 =>	x"27272727",
		582 =>	x"27272727",
		583 =>	x"27272727",
		584 =>	x"27272727",
		585 =>	x"27272727",
		586 =>	x"27272727",
		587 =>	x"27272727",
		588 =>	x"27272727",
		589 =>	x"27272727",
		590 =>	x"27272727",
		591 =>	x"27272727",
		592 =>	x"27272727",
		593 =>	x"27272727",
		594 =>	x"27272727",
		595 =>	x"27272727",
		596 =>	x"27272727",
		597 =>	x"27272727",
		598 =>	x"27272727",
		599 =>	x"27272727",
		600 =>	x"27272727",
		601 =>	x"27272727",
		602 =>	x"27272727",
		603 =>	x"27272727",
		604 =>	x"27272727",
		605 =>	x"27272727",
		606 =>	x"27272727",
		607 =>	x"27272727",
		608 =>	x"27272727",
		609 =>	x"27272727",
		610 =>	x"27272727",
		611 =>	x"27272727",
		612 =>	x"27272727",
		613 =>	x"27272727",
		614 =>	x"27272727",
		615 =>	x"27272727",
		616 =>	x"27272727",
		617 =>	x"27272727",
		618 =>	x"27272727",
		619 =>	x"27272727",
		620 =>	x"27272727",
		621 =>	x"27272727",
		622 =>	x"27272727",
		623 =>	x"27272727",
		624 =>	x"27272727",
		625 =>	x"27272727",
		626 =>	x"27272727",
		627 =>	x"27272727",
		628 =>	x"27272727",
		629 =>	x"27272727",
		630 =>	x"27272727",
		631 =>	x"27272727",
		632 =>	x"27272727",
		633 =>	x"27272727",
		634 =>	x"27272727",
		635 =>	x"27272727",
		636 =>	x"27272727",
		637 =>	x"27272727",
		638 =>	x"27272727",
		639 =>	x"1F1C2008", -- IMG_16x18_tobla3
		640 =>	x"080B250B",
		641 =>	x"0B252508",
		642 =>	x"08081C1F",
		643 =>	x"1C1C0808",
		644 =>	x"25090925",
		645 =>	x"09092508",
		646 =>	x"08081C1C",
		647 =>	x"1C080808",
		648 =>	x"25250925",
		649 =>	x"0A250808",
		650 =>	x"0B08081C",
		651 =>	x"1C080825",
		652 =>	x"250B2525",
		653 =>	x"25090925",
		654 =>	x"08081C1C",
		655 =>	x"1C1C0825",
		656 =>	x"25252509",
		657 =>	x"09090B08",
		658 =>	x"250B1C1E",
		659 =>	x"1C080825",
		660 =>	x"2525090D",
		661 =>	x"09092508",
		662 =>	x"2508081C",
		663 =>	x"1C08080B",
		664 =>	x"0B25090A",
		665 =>	x"0D0A0B08",
		666 =>	x"25081C1C",
		667 =>	x"1C08080B",
		668 =>	x"25090A09",
		669 =>	x"09090925",
		670 =>	x"09080808",
		671 =>	x"080B2525",
		672 =>	x"25090A09",
		673 =>	x"09090925",
		674 =>	x"2508081C",
		675 =>	x"1C080B25",
		676 =>	x"09090A09",
		677 =>	x"0A090925",
		678 =>	x"090B081E",
		679 =>	x"1C080B25",
		680 =>	x"09090909",
		681 =>	x"09252509",
		682 =>	x"25080820",
		683 =>	x"1C080825",
		684 =>	x"09250909",
		685 =>	x"09250825",
		686 =>	x"25080808",
		687 =>	x"1E1C0825",
		688 =>	x"25250909",
		689 =>	x"2509250B",
		690 =>	x"081C1C1C",
		691 =>	x"1E1C080B",
		692 =>	x"25090925",
		693 =>	x"250B0808",
		694 =>	x"08081C1F",
		695 =>	x"1E1C2008",
		696 =>	x"25090925",
		697 =>	x"0B080808",
		698 =>	x"081C1C1E",
		699 =>	x"1F1E1C08",
		700 =>	x"0B090A25",
		701 =>	x"2525081C",
		702 =>	x"081C1C1E",



--			***** MAP *****


		703 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		704 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		705 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		706 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		707 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		708 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		709 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		710 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		711 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		712 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		713 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		714 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		715 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		716 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		717 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		718 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		719 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		720 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		721 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		722 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		723 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		724 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		725 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		726 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		727 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		728 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		729 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		730 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		731 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		732 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		733 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		734 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		735 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		736 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		737 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		738 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		739 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		740 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		741 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		742 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		743 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		744 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		745 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		746 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		747 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		748 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		749 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		750 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		751 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		752 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		753 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		754 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		755 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		756 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		757 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		758 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		759 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		760 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		761 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		762 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		763 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		764 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		765 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		766 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		767 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		768 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		769 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		770 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		771 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		772 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		773 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		774 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		775 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		776 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		777 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		778 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		779 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		780 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		781 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		782 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		783 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		784 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		785 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		786 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		787 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		788 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		789 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		790 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		791 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		792 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		793 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		794 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		795 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		796 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		797 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		798 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		799 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		800 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		801 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		802 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		803 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		804 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		805 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		806 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		807 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		808 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		809 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		810 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		811 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		812 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		813 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		814 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		815 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		816 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		817 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		818 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		819 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		820 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		821 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		822 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		823 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		824 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		825 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		826 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		827 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		828 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		829 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		830 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		831 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		832 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		833 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		834 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		835 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		836 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		837 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		838 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		839 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		840 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		841 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		842 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		843 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		844 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		845 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		846 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		847 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		848 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		849 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		850 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		851 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		852 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		853 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		854 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		855 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		856 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		857 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		858 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		859 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		860 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		861 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		862 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		863 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		864 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		865 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		866 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		867 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		868 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		869 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		870 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		871 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		872 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		873 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		874 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		875 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		876 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		877 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		878 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		879 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		880 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		881 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		882 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		883 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		884 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		885 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		886 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		887 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		888 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		889 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		890 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		891 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		892 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		893 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		894 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		895 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		896 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		897 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		898 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		899 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		900 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		901 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		902 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		903 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		904 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		905 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		906 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		907 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		908 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		909 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		910 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		911 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		912 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		913 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		914 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		915 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		916 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		917 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		918 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		919 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		920 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		921 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		922 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		923 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		924 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		925 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		926 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		927 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		928 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		929 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		930 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		931 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		932 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		933 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		934 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		935 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		936 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		937 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		938 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		939 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		940 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		941 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		942 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		943 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		944 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		945 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		946 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		947 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		948 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		949 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		950 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		951 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		952 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		953 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		954 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		955 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		956 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		957 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		958 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		959 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		960 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		961 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		962 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		963 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		964 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		965 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		966 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		967 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		968 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		969 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		970 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		971 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		972 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		973 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		974 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		975 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		976 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		977 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		978 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		979 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		980 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		981 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		982 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		983 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		984 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		985 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		986 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		987 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		988 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		989 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		990 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		991 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		992 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		993 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		994 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		995 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		996 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		997 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		998 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		999 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1000 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1001 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1002 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1003 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1004 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1005 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1006 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1007 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1008 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1009 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1010 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1011 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1012 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1013 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1014 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1015 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1016 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1017 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1018 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1019 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1020 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1021 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1022 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1023 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1024 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1025 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1026 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1027 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1028 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1029 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1030 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1031 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1032 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1033 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1034 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1035 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1036 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1037 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1038 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1039 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1040 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1041 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1042 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1043 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1044 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1045 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1046 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1047 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1048 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1049 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1050 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1051 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1052 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1053 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1054 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1055 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1056 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1057 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1058 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1059 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1060 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1061 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1062 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1063 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1064 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1065 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1066 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1067 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1068 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1069 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1070 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1071 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1072 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1073 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1074 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1075 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1076 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1077 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1078 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1079 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1080 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1081 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1082 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1083 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1084 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1085 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1086 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1087 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1088 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1089 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1090 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1091 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1092 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1093 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1094 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1095 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1096 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1097 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1098 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1099 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1100 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1101 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1102 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1103 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1104 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1105 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1106 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1107 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1108 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1109 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1110 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1111 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1112 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1113 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1114 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1115 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1116 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1117 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1118 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1119 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1120 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1121 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1122 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1123 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1124 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1125 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1126 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1127 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1128 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1129 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1130 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1131 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1132 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1133 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1134 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1135 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1136 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1137 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1138 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1139 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1140 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1141 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1142 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1143 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1144 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1145 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1146 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1147 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1148 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1149 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1150 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1151 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1152 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1153 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1154 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1155 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1156 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1157 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1158 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1159 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1160 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1161 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1162 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1163 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1164 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1165 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1166 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1167 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1168 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1169 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1170 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1171 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1172 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1173 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1174 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1175 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1176 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1177 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1178 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1179 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1180 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1181 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1182 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1183 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1184 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1185 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1186 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1187 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1188 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1189 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1190 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1191 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1192 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1193 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1194 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1195 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1196 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1197 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1198 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1199 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1200 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1201 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1202 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1203 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1204 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1205 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1206 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1207 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1208 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1209 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1210 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1211 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1212 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1213 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1214 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1215 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1216 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1217 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1218 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1219 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1220 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1221 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1222 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1223 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1224 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1225 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1226 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1227 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1228 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1229 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1230 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1231 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1232 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1233 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1234 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1235 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1236 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1237 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1238 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1239 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1240 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1241 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1242 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1243 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1244 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1245 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1246 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1247 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1248 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1249 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1250 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1251 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1252 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1253 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1254 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1255 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1256 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1257 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1258 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1259 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1260 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1261 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1262 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1263 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1264 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1265 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1266 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1267 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1268 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1269 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1270 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1271 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1272 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1273 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1274 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1275 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1276 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1277 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1278 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1279 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1280 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1281 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1282 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1283 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1284 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1285 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1286 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1287 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1288 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1289 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1290 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1291 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1292 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1293 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1294 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1295 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1296 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1297 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1298 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1299 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1300 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1301 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1302 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1303 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1304 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1305 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1306 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1307 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1308 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1309 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1310 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1311 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1312 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1313 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1314 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1315 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1316 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1317 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1318 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1319 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1320 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1321 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1322 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1323 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1324 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1325 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1326 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1327 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1328 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1329 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1330 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1331 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1332 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1333 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1334 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1335 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1336 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1337 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1338 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1339 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1340 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1341 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1342 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1343 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1344 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1345 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1346 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1347 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1348 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1349 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1350 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1351 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1352 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1353 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1354 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1355 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1356 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1357 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1358 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1359 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1360 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1361 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1362 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1363 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1364 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1365 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1366 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1367 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1368 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1369 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1370 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1371 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1372 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1373 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1374 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1375 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1376 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1377 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1378 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1379 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1380 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1381 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1382 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1383 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1384 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1385 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1386 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1387 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1388 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1389 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1390 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1391 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1392 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1393 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1394 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1395 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1396 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1397 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1398 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1399 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1400 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1401 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1402 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1403 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1404 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1405 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1406 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1407 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1408 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1409 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1410 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1411 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1412 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1413 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1414 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1415 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1416 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1417 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1418 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1419 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1420 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1421 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1422 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1423 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1424 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1425 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1426 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1427 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1428 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1429 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1430 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1431 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1432 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1433 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1434 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1435 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1436 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1437 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1438 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1439 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1440 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1441 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1442 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1443 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1444 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1445 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1446 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1447 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1448 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1449 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1450 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1451 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1452 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1453 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1454 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1455 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1456 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1457 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1458 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1459 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1460 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1461 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1462 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1463 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1464 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1465 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1466 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1467 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1468 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1469 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1470 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1471 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1472 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1473 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1474 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1475 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1476 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1477 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1478 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1479 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1480 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1481 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1482 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1483 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1484 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1485 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1486 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1487 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1488 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1489 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1490 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1491 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1492 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1493 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1494 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1495 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1496 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1497 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1498 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1499 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1500 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1501 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1502 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1503 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1504 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1505 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1506 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1507 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1508 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1509 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1510 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1511 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1512 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1513 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1514 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1515 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1516 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1517 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1518 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1519 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1520 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1521 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1522 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1523 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1524 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1525 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1526 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1527 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1528 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1529 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1530 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1531 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1532 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1533 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1534 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1535 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1536 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1537 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1538 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1539 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1540 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1541 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1542 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1543 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1544 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1545 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1546 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1547 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1548 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1549 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1550 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1551 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1552 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1553 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1554 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1555 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1556 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1557 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1558 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1559 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1560 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1561 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1562 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1563 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1564 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1565 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1566 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1567 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1568 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1569 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1570 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1571 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1572 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1573 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1574 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1575 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1576 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1577 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1578 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1579 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1580 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1581 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1582 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1583 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1584 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1585 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1586 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1587 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1588 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1589 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1590 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1591 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1592 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1593 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1594 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1595 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1596 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1597 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1598 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1599 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1600 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1601 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1602 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1603 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1604 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1605 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1606 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1607 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1608 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1609 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1610 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1611 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1612 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1613 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1614 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1615 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1616 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1617 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1618 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1619 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1620 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1621 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1622 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1623 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1624 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1625 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1626 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1627 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1628 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1629 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1630 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1631 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1632 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1633 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1634 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1635 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1636 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1637 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1638 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1639 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1640 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1641 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1642 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1643 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1644 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1645 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1646 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1647 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1648 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1649 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1650 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1651 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1652 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1653 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1654 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1655 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1656 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1657 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1658 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1659 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1660 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1661 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1662 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1663 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1664 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1665 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1666 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1667 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1668 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1669 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1670 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1671 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1672 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1673 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1674 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1675 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1676 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1677 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1678 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1679 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1680 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1681 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1682 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1683 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1684 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1685 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1686 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1687 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1688 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1689 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1690 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1691 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1692 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1693 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1694 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1695 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1696 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1697 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1698 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1699 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1700 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1701 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1702 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1703 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1704 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1705 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1706 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1707 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1708 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1709 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1710 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1711 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1712 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1713 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1714 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1715 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1716 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1717 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1718 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1719 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1720 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1721 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1722 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1723 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1724 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1725 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1726 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1727 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1728 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1729 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1730 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1731 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1732 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1733 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1734 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1735 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1736 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1737 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1738 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1739 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1740 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1741 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1742 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1743 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1744 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1745 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1746 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1747 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1748 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1749 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1750 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1751 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1752 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1753 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1754 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1755 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1756 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1757 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1758 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1759 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1760 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1761 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1762 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1763 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1764 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1765 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1766 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1767 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1768 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1769 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1770 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1771 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1772 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1773 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1774 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1775 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1776 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1777 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1778 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1779 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1780 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1781 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1782 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1783 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1784 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1785 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1786 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1787 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1788 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1789 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1790 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1791 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1792 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1793 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1794 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1795 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1796 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1797 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1798 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1799 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1800 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1801 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1802 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1803 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1804 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1805 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1806 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1807 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1808 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1809 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1810 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1811 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1812 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1813 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1814 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1815 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1816 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1817 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1818 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1819 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1820 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1821 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1822 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1823 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1824 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1825 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1826 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1827 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1828 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1829 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1830 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1831 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1832 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1833 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1834 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1835 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1836 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1837 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1838 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1839 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1840 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1841 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1842 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1843 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1844 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1845 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1846 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1847 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1848 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1849 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1850 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1851 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1852 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1853 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1854 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1855 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1856 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1857 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1858 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1859 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1860 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1861 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1862 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1863 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1864 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1865 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1866 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1867 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1868 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1869 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1870 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1871 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1872 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1873 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1874 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1875 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1876 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1877 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1878 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1879 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1880 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1881 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1882 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1883 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1884 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1885 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1886 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1887 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1888 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1889 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1890 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1891 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1892 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1893 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1894 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1895 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1896 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1897 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1898 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1899 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1900 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1901 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1902 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		others => x"00000000"
	);


begin

	process(i_clk)
	begin
		if rising_edge(i_clk) then
			-- memory write --
			if i_we = '1' then
				mem(to_integer(unsigned(i_w_addr))) <= i_data;
			end if;
			-- memory read -- 
			o_data <= mem(to_integer(unsigned(i_r_addr)));
			
		end if; 
	end process;

end architecture arch;

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity ram is
	generic
	(
		DATA_WIDTH : natural := 32;		    -- 4 byte one line of memory
		ADDR_WIDTH : natural := 13			    -- 24576 bytes size of memory
	);

	port(
		i_clk    : in  std_logic;
		i_r_addr : in  std_logic_vector(ADDR_WIDTH-1 downto 0);
		i_data   : in  std_logic_vector(DATA_WIDTH-1 downto 0);
		i_we     : in  std_logic;
		i_w_addr : in  std_logic_vector(ADDR_WIDTH-1 downto 0);
		o_data   : out std_logic_vector(DATA_WIDTH-1 downto 0)
	);
end entity ram;

architecture arch of ram is

	type ram_t is array (0 to 2**ADDR_WIDTH-1) of std_logic_vector(DATA_WIDTH-1 downto 0);


-- GENERATED BY BC_MEM_PACKER

-- DATE: Thu May 18 16:01:02 2017

	signal mem : ram_t := (

--			***** COLOR PALLETE *****



		0 =>	x"00000000", -- R: 0 G: 0 B: 0
		1 =>	x"00004009", -- R: 9 G: 64 B: 0
		2 =>	x"00001E74", -- R: 116 G: 30 B: 0
		3 =>	x"00FC7F22", -- R: 34 G: 127 B: 252
		4 =>	x"00710008", -- R: 8 G: 0 B: 113
		5 =>	x"00800000", -- R: 0 G: 0 B: 128
		6 =>	x"00000400", -- R: 0 G: 4 B: 0
		7 =>	x"00010000", -- R: 0 G: 0 B: 1
		8 =>	x"00F8A659", -- R: 89 G: 166 B: 248
		9 =>	x"0000B108", -- R: 8 G: 177 B: 0
		10 =>	x"00000009", -- R: 9 G: 0 B: 0
		11 =>	x"00040100", -- R: 0 G: 1 B: 4
		12 =>	x"00001200", -- R: 0 G: 18 B: 0
		13 =>	x"00001252", -- R: 82 G: 18 B: 0
		14 =>	x"00710000", -- R: 0 G: 0 B: 113
		15 =>	x"0000AC59", -- R: 89 G: 172 B: 0
		16 =>	x"0000C8DE", -- R: 222 G: 200 B: 0
		17 =>	x"00590000", -- R: 0 G: 0 B: 89
		18 =>	x"00FFFFFF", -- R: 255 G: 255 B: 255
		19 =>	x"00FFFFF6", -- R: 246 G: 255 B: 255
		20 =>	x"0007FFFF", -- R: 255 G: 255 B: 7
		21 =>	x"00FFFDFD", -- R: 253 G: 253 B: 255
		22 =>	x"00FDFD00", -- R: 0 G: 253 B: 253
		23 =>	x"003A74FD", -- R: 253 G: 116 B: 58
		24 =>	x"005A3171", -- R: 113 G: 49 B: 90
		25 =>	x"00AC5900", -- R: 0 G: 89 B: 172
		26 =>	x"00788655", -- R: 85 G: 134 B: 120
		27 =>	x"00FF07A6", -- R: 166 G: 7 B: 255
		28 =>	x"005DAFAF", -- R: 175 G: 175 B: 93
		29 =>	x"00AEF6FF", -- R: 255 G: 246 B: 174
		30 =>	x"00A400AD", -- R: 173 G: 0 B: 164
		31 =>	x"005CA5FF", -- R: 255 G: 165 B: 92
		32 =>	x"00FFF608", -- R: 8 G: 246 B: 255
		33 =>	x"00FF5252", -- R: 82 G: 82 B: 255
		34 =>	x"00A69FA7", -- R: 167 G: 159 B: 166
		35 =>	x"000707AF", -- R: 175 G: 7 B: 7
		36 =>	x"000707FF", -- R: 255 G: 7 B: 7
		37 =>	x"0008A4F6", -- R: 246 G: 164 B: 8
		38 =>	x"00FF9EA7", -- R: 167 G: 158 B: 255
		39 =>	x"00A7AFAF", -- R: 175 G: 175 B: 167
		40 =>	x"00A7AF07", -- R: 7 G: 175 B: 167
		41 =>	x"00FFFFAE", -- R: 174 G: 255 B: 255
		42 =>	x"00AFAFAF", -- R: 175 G: 175 B: 175
		43 =>	x"00FFF607", -- R: 7 G: 246 B: 255
		44 =>	x"000707A4", -- R: 164 G: 7 B: 7
		45 =>	x"0099A3A3", -- R: 163 G: 163 B: 153
		46 =>	x"005B1453", -- R: 83 G: 20 B: 91
		47 =>	x"00A3A3F7", -- R: 247 G: 163 B: 163
		48 =>	x"009EA5F7", -- R: 247 G: 165 B: 158
		49 =>	x"00F7F7F7", -- R: 247 G: 247 B: 247
		50 =>	x"00ECEBA3", -- R: 163 G: 235 B: 236
		51 =>	x"009AA4FF", -- R: 255 G: 164 B: 154
		52 =>	x"00FFFF07", -- R: 7 G: 255 B: 255
		53 =>	x"009EA7AF", -- R: 175 G: 167 B: 158
		54 =>	x"00B7AFAF", -- R: 175 G: 175 B: 183
		55 =>	x"00F708A4", -- R: 164 G: 8 B: 247
		56 =>	x"00A39BAC", -- R: 172 G: 155 B: 163
		57 =>	x"00F65B0A", -- R: 10 G: 91 B: 246
		58 =>	x"000A549F", -- R: 159 G: 84 B: 10
		59 =>	x"009FA7AF", -- R: 175 G: 167 B: 159
		60 =>	x"00A7A607", -- R: 7 G: 166 B: 167
		61 =>	x"00FFF65C", -- R: 92 G: 246 B: 255
		62 =>	x"0014130A", -- R: 10 G: 19 B: 20
		63 =>	x"0054A6A5", -- R: 165 G: 166 B: 84
		64 =>	x"00535E9E", -- R: 158 G: 94 B: 83
		65 =>	x"00A607FF", -- R: 255 G: 7 B: 166
		66 =>	x"005C141C", -- R: 28 G: 20 B: 92
		67 =>	x"0014A3EC", -- R: 236 G: 163 B: 20
		68 =>	x"00EC9A13", -- R: 19 G: 154 B: 236
		69 =>	x"00145C5B", -- R: 91 G: 92 B: 20
		70 =>	x"00F7F6FF", -- R: 255 G: 246 B: 247
		71 =>	x"0008F6F6", -- R: 246 G: 246 B: 8
		72 =>	x"000808F6", -- R: 246 G: 8 B: 8
		73 =>	x"00F6F6FF", -- R: 255 G: 246 B: 246
		74 =>	x"00FFFFF7", -- R: 247 G: 255 B: 255
		75 =>	x"005B0A5C", -- R: 92 G: 10 B: 91
		76 =>	x"009E9E5D", -- R: 93 G: 158 B: 158
		77 =>	x"00A6AFAE", -- R: 174 G: 175 B: 166
		78 =>	x"0007F6FF", -- R: 255 G: 246 B: 7
		79 =>	x"00AEAFAF", -- R: 175 G: 175 B: 174
		80 =>	x"005DA607", -- R: 7 G: 166 B: 93
		81 =>	x"00FFA55C", -- R: 92 G: 165 B: 255
		82 =>	x"00AD00A4", -- R: 164 G: 0 B: 173
		83 =>	x"00FFFF52", -- R: 82 G: 255 B: 255
		84 =>	x"0052FF08", -- R: 8 G: 255 B: 82
		85 =>	x"00F6FFFF", -- R: 255 G: 255 B: 246
		86 =>	x"00FFF6A4", -- R: 164 G: 246 B: 255
		87 =>	x"0008FF07", -- R: 7 G: 255 B: 8
		88 =>	x"0007AF07", -- R: 7 G: 175 B: 7
		89 =>	x"0007A79F", -- R: 159 G: 167 B: 7
		90 =>	x"00A6FFFF", -- R: 255 G: 255 B: 166
		91 =>	x"0007AFA7", -- R: 167 G: 175 B: 7
		92 =>	x"00AFAFA7", -- R: 167 G: 175 B: 175
		93 =>	x"00A79EFF", -- R: 255 G: 158 B: 167
		94 =>	x"00FF07AF", -- R: 175 G: 7 B: 255
		95 =>	x"00AFA7AE", -- R: 174 G: 167 B: 175
		96 =>	x"00FFF7A3", -- R: 163 G: 247 B: 255
		97 =>	x"00A35314", -- R: 20 G: 83 B: 163
		98 =>	x"005BA3A3", -- R: 163 G: 163 B: 91
		99 =>	x"0099A407", -- R: 7 G: 164 B: 153
		100 =>	x"000707F6", -- R: 246 G: 7 B: 7
		101 =>	x"00FFA49A", -- R: 154 G: 164 B: 255
		102 =>	x"00A3EBEC", -- R: 236 G: 235 B: 163
		103 =>	x"00F7A59E", -- R: 158 G: 165 B: 247
		104 =>	x"00AEFFFF", -- R: 255 G: 255 B: 174
		105 =>	x"00FFFFAC", -- R: 172 G: 255 B: 255
		106 =>	x"009BA3A4", -- R: 164 G: 163 B: 155
		107 =>	x"0008F7AF", -- R: 175 G: 247 B: 8
		108 =>	x"00AFB7AF", -- R: 175 G: 183 B: 175
		109 =>	x"00A79E07", -- R: 7 G: 158 B: 167
		110 =>	x"00A7AFA7", -- R: 167 G: 175 B: 167
		111 =>	x"009F9F54", -- R: 84 G: 159 B: 159
		112 =>	x"000A0A5B", -- R: 91 G: 10 B: 10
		113 =>	x"009E5E53", -- R: 83 G: 94 B: 158
		114 =>	x"00A5A654", -- R: 84 G: 166 B: 165
		115 =>	x"000A1314", -- R: 20 G: 19 B: 10
		116 =>	x"005CF6FF", -- R: 255 G: 246 B: 92
		117 =>	x"00F6F75B", -- R: 91 G: 247 B: 246
		118 =>	x"005C1413", -- R: 19 G: 20 B: 92
		119 =>	x"009AECEC", -- R: 236 G: 236 B: 154
		120 =>	x"00A3141C", -- R: 28 G: 20 B: 163
		121 =>	x"00145CFF", -- R: 255 G: 92 B: 20
		122 =>	x"00FFF6F6", -- R: 246 G: 246 B: 255
		123 =>	x"00F60808", -- R: 8 G: 8 B: 246
		124 =>	x"00F6F608", -- R: 8 G: 246 B: 246
		125 =>	x"00F6AEAE", -- R: 174 G: 174 B: 246
		126 =>	x"00AFA65D", -- R: 93 G: 166 B: 175
		127 =>	x"009E9E5C", -- R: 92 G: 158 B: 158
		128 =>	x"000A5BF7", -- R: 247 G: 91 B: 10
		129 =>	x"00E8E8E8", -- R: 232 G: 232 B: 232
		130 =>	x"00E8FDFD", -- R: 253 G: 253 B: 232
		131 =>	x"005D5D5C", -- R: 92 G: 93 B: 93
		132 =>	x"005C545D", -- R: 93 G: 84 B: 92
		133 =>	x"00545C5D", -- R: 93 G: 92 B: 84
		134 =>	x"005D5454", -- R: 84 G: 84 B: 93
		135 =>	x"0054545D", -- R: 93 G: 84 B: 84
		136 =>	x"005DFDFD", -- R: 253 G: 253 B: 93
		137 =>	x"005C5D5C", -- R: 92 G: 93 B: 92
		138 =>	x"005D5D5D", -- R: 93 G: 93 B: 93
		139 =>	x"00545C5C", -- R: 92 G: 92 B: 84
		140 =>	x"00545454", -- R: 84 G: 84 B: 84
		141 =>	x"005D545D", -- R: 93 G: 84 B: 93
		142 =>	x"009D5C5D", -- R: 93 G: 92 B: 157
		143 =>	x"005C549D", -- R: 157 G: 84 B: 92
		144 =>	x"005D549D", -- R: 157 G: 84 B: 93
		145 =>	x"005C5D5D", -- R: 93 G: 93 B: 92
		146 =>	x"005C9D5D", -- R: 93 G: 157 B: 92
		147 =>	x"00A55C5C", -- R: 92 G: 92 B: 165
		148 =>	x"005D5DA5", -- R: 165 G: 93 B: 93
		149 =>	x"005C54A5", -- R: 165 G: 84 B: 92
		150 =>	x"005D5C5D", -- R: 93 G: 92 B: 93
		151 =>	x"005D5C5C", -- R: 92 G: 92 B: 93
		152 =>	x"005D9D5C", -- R: 92 G: 157 B: 93
		153 =>	x"005D540B", -- R: 11 G: 84 B: 93
		154 =>	x"005D9D5D", -- R: 93 G: 157 B: 93
		155 =>	x"00A6A5A6", -- R: 166 G: 165 B: 166
		156 =>	x"00A55D5D", -- R: 93 G: 93 B: 165
		157 =>	x"005D5C9D", -- R: 157 G: 92 B: 93
		158 =>	x"005D5D9D", -- R: 157 G: 93 B: 93
		159 =>	x"00A6A55D", -- R: 93 G: 165 B: 166
		160 =>	x"005CA65D", -- R: 93 G: 166 B: 92
		161 =>	x"00A6545C", -- R: 92 G: 84 B: 166
		162 =>	x"009D5D5D", -- R: 93 G: 93 B: 157
		163 =>	x"00A65D5D", -- R: 93 G: 93 B: 166
		164 =>	x"005D5D54", -- R: 84 G: 93 B: 93
		165 =>	x"00A6545D", -- R: 93 G: 84 B: 166
		166 =>	x"005D54A6", -- R: 166 G: 84 B: 93
		167 =>	x"005DA654", -- R: 84 G: 166 B: 93
		168 =>	x"005C5D9D", -- R: 157 G: 93 B: 92
		169 =>	x"00545D5D", -- R: 93 G: 93 B: 84
		170 =>	x"005D655D", -- R: 93 G: 101 B: 93
		171 =>	x"005D5DA6", -- R: 166 G: 93 B: 93
		172 =>	x"00545D54", -- R: 84 G: 93 B: 84
		173 =>	x"005DA69D", -- R: 157 G: 166 B: 93
		174 =>	x"00545DA6", -- R: 166 G: 93 B: 84
		175 =>	x"005DA65D", -- R: 93 G: 166 B: 93
		176 =>	x"00A65D9D", -- R: 157 G: 93 B: 166
		177 =>	x"005D0B5D", -- R: 93 G: 11 B: 93
		178 =>	x"005D4B54", -- R: 84 G: 75 B: 93
		179 =>	x"00545D5C", -- R: 92 G: 93 B: 84
		180 =>	x"00666666", -- R: 102 G: 102 B: 102
		181 =>	x"0066FDFD", -- R: 253 G: 253 B: 102
		182 =>	x"000A5354", -- R: 84 G: 83 B: 10
		183 =>	x"005C5C5D", -- R: 93 G: 92 B: 92
		184 =>	x"00655D5D", -- R: 93 G: 93 B: 101
		185 =>	x"0065655C", -- R: 92 G: 101 B: 101
		186 =>	x"005C5C53", -- R: 83 G: 92 B: 92
		187 =>	x"000AFDFD", -- R: 253 G: 253 B: 10
		188 =>	x"00535C5C", -- R: 92 G: 92 B: 83
		189 =>	x"0065655D", -- R: 93 G: 101 B: 101
		190 =>	x"00656565", -- R: 101 G: 101 B: 101
		191 =>	x"00A5A565", -- R: 101 G: 165 B: 165
		192 =>	x"0053535C", -- R: 92 G: 83 B: 83
		193 =>	x"005C5C65", -- R: 101 G: 92 B: 92
		194 =>	x"0065A565", -- R: 101 G: 165 B: 101
		195 =>	x"00A6655C", -- R: 92 G: 101 B: 166
		196 =>	x"005C5353", -- R: 83 G: 83 B: 92
		197 =>	x"0065A5A5", -- R: 165 G: 165 B: 101
		198 =>	x"00655C5C", -- R: 92 G: 92 B: 101
		199 =>	x"005D5D65", -- R: 101 G: 93 B: 93
		200 =>	x"00A5A6AE", -- R: 174 G: 166 B: 165
		201 =>	x"00A65D5C", -- R: 92 G: 93 B: 166
		202 =>	x"00655C53", -- R: 83 G: 92 B: 101
		203 =>	x"005C6565", -- R: 101 G: 101 B: 92
		204 =>	x"0065A5AE", -- R: 174 G: 165 B: 101
		205 =>	x"005C655C", -- R: 92 G: 101 B: 92
		206 =>	x"00535C65", -- R: 101 G: 92 B: 83
		207 =>	x"00A5A5A5", -- R: 165 G: 165 B: 165
		208 =>	x"005D5C65", -- R: 101 G: 92 B: 93
		209 =>	x"005D5313", -- R: 19 G: 83 B: 93
		210 =>	x"00535C5D", -- R: 93 G: 92 B: 83
		211 =>	x"00A55D5C", -- R: 92 G: 93 B: 165
		212 =>	x"00135C5D", -- R: 93 G: 92 B: 19
		213 =>	x"00A5A6A5", -- R: 165 G: 166 B: 165
		214 =>	x"0065A5A6", -- R: 166 G: 165 B: 101
		215 =>	x"00A565A5", -- R: 165 G: 101 B: 165
		216 =>	x"005C5C5C", -- R: 92 G: 92 B: 92
		217 =>	x"0013535C", -- R: 92 G: 83 B: 19
		218 =>	x"00A5655D", -- R: 93 G: 101 B: 165
		219 =>	x"005C65A5", -- R: 165 G: 101 B: 92
		220 =>	x"00A5655C", -- R: 92 G: 101 B: 165
		221 =>	x"005C5D65", -- R: 101 G: 93 B: 92
		222 =>	x"005C5C54", -- R: 84 G: 92 B: 92
		223 =>	x"000A1353", -- R: 83 G: 19 B: 10
		224 =>	x"005C5DA5", -- R: 165 G: 93 B: 92
		225 =>	x"00A66565", -- R: 101 G: 101 B: 166
		226 =>	x"00131353", -- R: 83 G: 19 B: 19
		227 =>	x"00545C65", -- R: 101 G: 92 B: 84
		228 =>	x"00531313", -- R: 19 G: 19 B: 83
		229 =>	x"005C530A", -- R: 10 G: 83 B: 92
		230 =>	x"00000000", -- Unused
		231 =>	x"00000000", -- Unused
		232 =>	x"00000000", -- Unused
		233 =>	x"00000000", -- Unused
		234 =>	x"00000000", -- Unused
		235 =>	x"00000000", -- Unused
		236 =>	x"00000000", -- Unused
		237 =>	x"00000000", -- Unused
		238 =>	x"00000000", -- Unused
		239 =>	x"00000000", -- Unused
		240 =>	x"00000000", -- Unused
		241 =>	x"00000000", -- Unused
		242 =>	x"00000000", -- Unused
		243 =>	x"00000000", -- Unused
		244 =>	x"00000000", -- Unused
		245 =>	x"00000000", -- Unused
		246 =>	x"00000000", -- Unused
		247 =>	x"00000000", -- Unused
		248 =>	x"00000000", -- Unused
		249 =>	x"00000000", -- Unused
		250 =>	x"00000000", -- Unused
		251 =>	x"00000000", -- Unused
		252 =>	x"00000000", -- Unused
		253 =>	x"00000000", -- Unused
		254 =>	x"00000000", -- Unused
--			***** 16x16 IMAGES *****




		255 =>	x"01000000", -- IMG_16x18_crvcina_desno
		256 =>	x"00000000",
		257 =>	x"00000000",
		258 =>	x"00000000",
		259 =>	x"00000000",
		260 =>	x"00020304",
		261 =>	x"05060700",
		262 =>	x"08090A0B",
		263 =>	x"00000000",
		264 =>	x"00000000",
		265 =>	x"00000000",
		266 =>	x"00000000",
		267 =>	x"00000000",
		268 =>	x"00000000",
		269 =>	x"00000000",
		270 =>	x"00000000",
		271 =>	x"00000000",
		272 =>	x"000C0D0E",
		273 =>	x"0F101100",
		274 =>	x"00000000",
		275 =>	x"00000000",
		276 =>	x"00000000",
		277 =>	x"00000000",
		278 =>	x"00000000",
		279 =>	x"00000000",
		280 =>	x"00000000",
		281 =>	x"00000000",
		282 =>	x"00000000",
		283 =>	x"00000000",
		284 =>	x"00000000",
		285 =>	x"00000000",
		286 =>	x"00000000",
		287 =>	x"00000000",
		288 =>	x"00000000",
		289 =>	x"00000000",
		290 =>	x"00000000",
		291 =>	x"00000000",
		292 =>	x"00000000",
		293 =>	x"00000000",
		294 =>	x"00000000",
		295 =>	x"12121314",
		296 =>	x"12151600",
		297 =>	x"17180019",
		298 =>	x"1A000000",
		299 =>	x"121B1C1D",
		300 =>	x"1212121E",
		301 =>	x"1F121212",
		302 =>	x"20211212",
		303 =>	x"12222324",
		304 =>	x"25122627",
		305 =>	x"28121229",
		306 =>	x"272A1412",
		307 =>	x"2B2C2D2E",
		308 =>	x"2F122930",
		309 =>	x"31323334",
		310 =>	x"35363738",
		311 =>	x"393A3B3C",
		312 =>	x"123D3E3F",
		313 =>	x"40411242",
		314 =>	x"43444546",
		315 =>	x"12121212",
		316 =>	x"12134748",
		317 =>	x"49124A4B",
		318 =>	x"4C4D1D12",
		319 =>	x"01000000", -- IMG_16x18_crvcina_levo
		320 =>	x"00000000",
		321 =>	x"00000000",
		322 =>	x"00000000",
		323 =>	x"00000000",
		324 =>	x"00020304",
		325 =>	x"05060700",
		326 =>	x"08090A0B",
		327 =>	x"00000000",
		328 =>	x"00000000",
		329 =>	x"00000000",
		330 =>	x"00000000",
		331 =>	x"00000000",
		332 =>	x"00000000",
		333 =>	x"00000000",
		334 =>	x"00000000",
		335 =>	x"00000000",
		336 =>	x"000C0D0E",
		337 =>	x"0F101100",
		338 =>	x"00000000",
		339 =>	x"00000000",
		340 =>	x"00000000",
		341 =>	x"00000000",
		342 =>	x"00000000",
		343 =>	x"00000000",
		344 =>	x"00000000",
		345 =>	x"00000000",
		346 =>	x"00000000",
		347 =>	x"00000000",
		348 =>	x"00000000",
		349 =>	x"00000000",
		350 =>	x"00000000",
		351 =>	x"00000000",
		352 =>	x"00000000",
		353 =>	x"00000000",
		354 =>	x"00000000",
		355 =>	x"00000000",
		356 =>	x"00000000",
		357 =>	x"00000000",
		358 =>	x"00000000",
		359 =>	x"12124E12",
		360 =>	x"12151600",
		361 =>	x"17180019",
		362 =>	x"1A000000",
		363 =>	x"12134F50",
		364 =>	x"12121251",
		365 =>	x"52121212",
		366 =>	x"53545512",
		367 =>	x"56575859",
		368 =>	x"5A12125B",
		369 =>	x"5C5D1212",
		370 =>	x"5E2A5F12",
		371 =>	x"60616263",
		372 =>	x"64656631",
		373 =>	x"6768696A",
		374 =>	x"6B6C6D12",
		375 =>	x"121B6E6F",
		376 =>	x"70551B71",
		377 =>	x"72737475",
		378 =>	x"76777879",
		379 =>	x"12121212",
		380 =>	x"1212127A",
		381 =>	x"7B7C5512",
		382 =>	x"7D7E7F80",
		383 =>	x"01000000", -- IMG_16x18_nebo_svetlo
		384 =>	x"00000000",
		385 =>	x"00000000",
		386 =>	x"00000000",
		387 =>	x"00000000",
		388 =>	x"00020304",
		389 =>	x"05060700",
		390 =>	x"08090A0B",
		391 =>	x"00000000",
		392 =>	x"00000000",
		393 =>	x"00000000",
		394 =>	x"00000000",
		395 =>	x"00000000",
		396 =>	x"00000000",
		397 =>	x"00000000",
		398 =>	x"00000000",
		399 =>	x"00000000",
		400 =>	x"000C0D0E",
		401 =>	x"0F101100",
		402 =>	x"00000000",
		403 =>	x"00000000",
		404 =>	x"00000000",
		405 =>	x"00000000",
		406 =>	x"00000000",
		407 =>	x"00000000",
		408 =>	x"00000000",
		409 =>	x"00000000",
		410 =>	x"00000000",
		411 =>	x"00000000",
		412 =>	x"00000000",
		413 =>	x"00000000",
		414 =>	x"00000000",
		415 =>	x"00000000",
		416 =>	x"00000000",
		417 =>	x"00000000",
		418 =>	x"00000000",
		419 =>	x"00000000",
		420 =>	x"00000000",
		421 =>	x"00000000",
		422 =>	x"00000000",
		423 =>	x"81818181",
		424 =>	x"81821600",
		425 =>	x"17180019",
		426 =>	x"1A000000",
		427 =>	x"81818181",
		428 =>	x"81818181",
		429 =>	x"81818181",
		430 =>	x"81818181",
		431 =>	x"81818181",
		432 =>	x"81818181",
		433 =>	x"81818181",
		434 =>	x"81818181",
		435 =>	x"81818181",
		436 =>	x"81818181",
		437 =>	x"81818181",
		438 =>	x"81818181",
		439 =>	x"81818181",
		440 =>	x"81818181",
		441 =>	x"81818181",
		442 =>	x"81818181",
		443 =>	x"81818181",
		444 =>	x"81818181",
		445 =>	x"81818181",
		446 =>	x"81818181",
		447 =>	x"01000000", -- IMG_16x18_oblak
		448 =>	x"00000000",
		449 =>	x"00000000",
		450 =>	x"00000000",
		451 =>	x"00000000",
		452 =>	x"00020304",
		453 =>	x"05060700",
		454 =>	x"08090A0B",
		455 =>	x"00000000",
		456 =>	x"00000000",
		457 =>	x"00000000",
		458 =>	x"00000000",
		459 =>	x"00000000",
		460 =>	x"00000000",
		461 =>	x"00000000",
		462 =>	x"00000000",
		463 =>	x"00000000",
		464 =>	x"000C0D0E",
		465 =>	x"0F101100",
		466 =>	x"00000000",
		467 =>	x"00000000",
		468 =>	x"00000000",
		469 =>	x"00000000",
		470 =>	x"00000000",
		471 =>	x"00000000",
		472 =>	x"00000000",
		473 =>	x"00000000",
		474 =>	x"00000000",
		475 =>	x"00000000",
		476 =>	x"00000000",
		477 =>	x"00000000",
		478 =>	x"00000000",
		479 =>	x"00000000",
		480 =>	x"00000000",
		481 =>	x"00000000",
		482 =>	x"00000000",
		483 =>	x"00000000",
		484 =>	x"00000000",
		485 =>	x"00000000",
		486 =>	x"00000000",
		487 =>	x"12121212",
		488 =>	x"12151600",
		489 =>	x"17180019",
		490 =>	x"1A000000",
		491 =>	x"12121212",
		492 =>	x"12121212",
		493 =>	x"12121212",
		494 =>	x"12121212",
		495 =>	x"12121212",
		496 =>	x"12121212",
		497 =>	x"12121212",
		498 =>	x"12121212",
		499 =>	x"12121212",
		500 =>	x"12121212",
		501 =>	x"12121212",
		502 =>	x"12121212",
		503 =>	x"12121212",
		504 =>	x"12121212",
		505 =>	x"12121212",
		506 =>	x"12121212",
		507 =>	x"12121212",
		508 =>	x"12121212",
		509 =>	x"12121212",
		510 =>	x"12121212",
		511 =>	x"01000000", -- IMG_16x18_tobla1
		512 =>	x"00000000",
		513 =>	x"00000000",
		514 =>	x"00000000",
		515 =>	x"00000000",
		516 =>	x"00020304",
		517 =>	x"05060700",
		518 =>	x"08090A0B",
		519 =>	x"00000000",
		520 =>	x"00000000",
		521 =>	x"00000000",
		522 =>	x"00000000",
		523 =>	x"00000000",
		524 =>	x"00000000",
		525 =>	x"00000000",
		526 =>	x"00000000",
		527 =>	x"00000000",
		528 =>	x"000C0D0E",
		529 =>	x"0F101100",
		530 =>	x"00000000",
		531 =>	x"00000000",
		532 =>	x"00000000",
		533 =>	x"00000000",
		534 =>	x"00000000",
		535 =>	x"00000000",
		536 =>	x"00000000",
		537 =>	x"00000000",
		538 =>	x"00000000",
		539 =>	x"00000000",
		540 =>	x"00000000",
		541 =>	x"00000000",
		542 =>	x"00000000",
		543 =>	x"00000000",
		544 =>	x"00000000",
		545 =>	x"00000000",
		546 =>	x"00000000",
		547 =>	x"00000000",
		548 =>	x"00000000",
		549 =>	x"00000000",
		550 =>	x"00000000",
		551 =>	x"83848586",
		552 =>	x"87881600",
		553 =>	x"17180019",
		554 =>	x"1A000000",
		555 =>	x"898A8B8A",
		556 =>	x"8C8D8E8D",
		557 =>	x"868C8687",
		558 =>	x"8F878A8C",
		559 =>	x"9091928A",
		560 =>	x"93949596",
		561 =>	x"978A8E97",
		562 =>	x"988D8799",
		563 =>	x"849A9B9C",
		564 =>	x"9D9E849F",
		565 =>	x"A0A18AA2",
		566 =>	x"8AA38AA4",
		567 =>	x"A5A6A4A4",
		568 =>	x"A7A883A9",
		569 =>	x"AAAB87A9",
		570 =>	x"8A97AC8A",
		571 =>	x"ADAEABAF",
		572 =>	x"8384B08D",
		573 =>	x"B18AB2AB",
		574 =>	x"B38A9CA3",
		575 =>	x"01000000", -- IMG_16x18_tobla2
		576 =>	x"00000000",
		577 =>	x"00000000",
		578 =>	x"00000000",
		579 =>	x"00000000",
		580 =>	x"00020304",
		581 =>	x"05060700",
		582 =>	x"08090A0B",
		583 =>	x"00000000",
		584 =>	x"00000000",
		585 =>	x"00000000",
		586 =>	x"00000000",
		587 =>	x"00000000",
		588 =>	x"00000000",
		589 =>	x"00000000",
		590 =>	x"00000000",
		591 =>	x"00000000",
		592 =>	x"000C0D0E",
		593 =>	x"0F101100",
		594 =>	x"00000000",
		595 =>	x"00000000",
		596 =>	x"00000000",
		597 =>	x"00000000",
		598 =>	x"00000000",
		599 =>	x"00000000",
		600 =>	x"00000000",
		601 =>	x"00000000",
		602 =>	x"00000000",
		603 =>	x"00000000",
		604 =>	x"00000000",
		605 =>	x"00000000",
		606 =>	x"00000000",
		607 =>	x"00000000",
		608 =>	x"00000000",
		609 =>	x"00000000",
		610 =>	x"00000000",
		611 =>	x"00000000",
		612 =>	x"00000000",
		613 =>	x"00000000",
		614 =>	x"00000000",
		615 =>	x"B4B4B4B4",
		616 =>	x"B4B51600",
		617 =>	x"17180019",
		618 =>	x"1A000000",
		619 =>	x"B4B4B4B4",
		620 =>	x"B4B4B4B4",
		621 =>	x"B4B4B4B4",
		622 =>	x"B4B4B4B4",
		623 =>	x"B4B4B4B4",
		624 =>	x"B4B4B4B4",
		625 =>	x"B4B4B4B4",
		626 =>	x"B4B4B4B4",
		627 =>	x"B4B4B4B4",
		628 =>	x"B4B4B4B4",
		629 =>	x"B4B4B4B4",
		630 =>	x"B4B4B4B4",
		631 =>	x"B4B4B4B4",
		632 =>	x"B4B4B4B4",
		633 =>	x"B4B4B4B4",
		634 =>	x"B4B4B4B4",
		635 =>	x"B4B4B4B4",
		636 =>	x"B4B4B4B4",
		637 =>	x"B4B4B4B4",
		638 =>	x"B4B4B4B4",
		639 =>	x"01000000", -- IMG_16x18_tobla3
		640 =>	x"00000000",
		641 =>	x"00000000",
		642 =>	x"00000000",
		643 =>	x"00000000",
		644 =>	x"00020304",
		645 =>	x"05060700",
		646 =>	x"08090A0B",
		647 =>	x"00000000",
		648 =>	x"00000000",
		649 =>	x"00000000",
		650 =>	x"00000000",
		651 =>	x"00000000",
		652 =>	x"00000000",
		653 =>	x"00000000",
		654 =>	x"00000000",
		655 =>	x"00000000",
		656 =>	x"000C0D0E",
		657 =>	x"0F101100",
		658 =>	x"00000000",
		659 =>	x"00000000",
		660 =>	x"00000000",
		661 =>	x"00000000",
		662 =>	x"00000000",
		663 =>	x"00000000",
		664 =>	x"00000000",
		665 =>	x"00000000",
		666 =>	x"00000000",
		667 =>	x"00000000",
		668 =>	x"00000000",
		669 =>	x"00000000",
		670 =>	x"00000000",
		671 =>	x"00000000",
		672 =>	x"00000000",
		673 =>	x"00000000",
		674 =>	x"00000000",
		675 =>	x"00000000",
		676 =>	x"00000000",
		677 =>	x"00000000",
		678 =>	x"00000000",
		679 =>	x"B6B7B8B9",
		680 =>	x"BABB1600",
		681 =>	x"17180019",
		682 =>	x"1A000000",
		683 =>	x"BCBDBEBF",
		684 =>	x"BAC0C1C2",
		685 =>	x"C389C4BC",
		686 =>	x"C5C5C6C4",
		687 =>	x"BCC7C8C9",
		688 =>	x"CAC0CBCC",
		689 =>	x"BFCDC4CE",
		690 =>	x"BECFD0D1",
		691 =>	x"D2C59BBF",
		692 =>	x"D3D4BED5",
		693 =>	x"CFB9C4B7",
		694 =>	x"D6CFD7D8",
		695 =>	x"D9BEBFDA",
		696 =>	x"C4C0DBC5",
		697 =>	x"DCB9BADD",
		698 =>	x"CFBFC2DE",
		699 =>	x"DFE0E1CA",
		700 =>	x"C4E2E3BF",
		701 =>	x"97BAE4D2",
		702 =>	x"C5BDD8E5",


--			***** MAP *****


		703 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		704 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		705 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		706 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		707 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		708 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		709 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		710 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		711 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		712 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		713 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		714 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		715 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		716 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		717 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		718 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		719 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		720 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		721 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		722 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		723 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		724 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		725 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		726 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		727 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		728 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		729 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		730 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		731 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		732 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		733 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		734 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		735 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		736 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		737 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		738 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		739 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		740 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		741 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		742 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		743 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		744 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		745 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		746 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		747 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		748 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		749 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		750 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		751 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		752 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		753 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		754 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		755 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		756 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		757 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		758 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		759 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		760 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		761 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		762 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		763 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		764 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		765 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		766 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		767 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		768 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		769 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		770 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		771 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		772 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		773 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		774 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		775 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		776 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		777 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		778 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		779 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		780 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		781 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		782 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		783 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		784 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		785 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		786 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		787 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		788 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		789 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		790 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		791 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		792 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		793 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		794 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		795 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		796 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		797 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		798 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		799 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		800 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		801 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		802 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		803 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		804 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		805 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		806 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		807 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		808 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		809 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		810 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		811 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		812 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		813 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		814 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		815 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		816 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		817 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		818 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		819 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		820 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		821 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		822 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		823 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		824 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		825 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		826 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		827 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		828 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		829 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		830 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		831 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		832 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		833 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		834 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		835 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		836 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		837 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		838 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		839 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		840 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		841 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		842 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		843 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		844 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		845 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		846 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		847 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		848 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		849 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		850 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		851 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		852 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		853 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		854 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		855 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		856 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		857 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		858 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		859 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		860 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		861 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		862 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		863 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		864 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		865 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		866 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		867 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		868 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		869 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		870 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		871 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		872 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		873 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		874 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		875 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		876 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		877 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		878 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		879 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		880 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		881 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		882 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		883 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		884 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		885 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		886 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		887 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		888 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		889 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		890 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		891 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		892 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		893 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		894 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		895 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		896 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		897 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		898 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		899 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		900 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		901 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		902 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		903 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		904 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		905 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		906 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		907 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		908 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		909 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		910 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		911 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		912 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		913 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		914 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		915 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		916 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		917 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		918 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		919 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		920 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		921 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		922 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		923 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		924 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		925 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		926 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		927 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		928 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		929 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		930 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		931 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		932 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		933 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		934 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		935 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		936 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		937 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		938 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		939 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		940 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		941 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		942 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		943 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		944 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		945 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		946 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		947 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		948 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		949 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		950 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		951 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		952 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		953 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		954 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		955 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		956 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		957 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		958 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		959 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		960 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		961 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		962 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		963 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		964 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		965 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		966 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		967 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		968 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		969 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		970 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		971 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		972 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		973 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		974 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		975 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		976 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		977 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		978 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		979 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		980 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		981 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		982 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		983 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		984 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		985 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		986 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		987 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		988 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		989 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		990 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		991 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		992 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		993 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		994 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		995 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		996 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		997 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		998 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		999 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1000 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1001 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1002 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1003 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1004 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1005 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1006 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1007 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1008 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1009 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1010 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1011 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1012 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1013 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1014 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1015 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1016 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1017 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1018 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1019 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1020 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1021 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1022 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1023 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1024 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1025 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1026 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1027 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1028 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1029 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1030 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1031 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1032 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1033 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1034 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1035 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1036 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1037 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1038 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1039 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1040 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1041 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1042 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1043 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1044 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1045 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1046 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1047 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1048 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1049 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1050 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1051 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1052 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1053 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1054 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1055 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1056 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1057 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1058 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1059 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1060 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1061 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1062 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1063 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1064 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1065 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1066 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1067 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1068 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1069 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1070 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1071 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1072 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1073 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1074 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1075 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1076 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1077 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1078 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1079 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1080 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1081 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1082 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1083 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1084 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1085 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1086 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1087 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1088 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1089 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1090 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1091 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1092 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1093 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1094 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1095 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1096 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1097 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1098 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1099 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1100 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1101 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1102 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1103 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1104 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1105 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1106 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1107 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1108 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1109 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1110 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1111 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1112 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1113 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1114 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1115 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1116 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1117 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1118 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1119 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1120 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1121 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1122 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1123 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1124 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1125 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1126 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1127 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1128 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1129 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1130 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1131 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1132 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1133 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1134 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1135 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1136 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1137 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1138 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1139 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1140 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1141 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1142 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1143 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1144 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1145 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1146 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1147 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1148 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1149 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1150 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1151 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1152 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1153 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1154 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1155 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1156 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1157 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1158 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1159 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1160 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1161 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1162 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1163 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1164 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1165 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1166 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1167 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1168 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1169 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1170 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1171 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1172 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1173 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1174 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1175 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1176 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1177 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1178 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1179 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1180 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1181 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1182 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1183 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1184 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1185 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1186 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1187 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1188 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1189 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1190 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1191 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1192 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1193 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1194 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1195 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1196 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1197 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1198 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1199 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1200 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1201 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1202 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1203 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1204 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1205 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1206 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1207 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1208 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1209 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1210 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1211 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1212 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1213 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1214 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1215 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1216 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1217 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1218 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1219 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1220 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1221 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1222 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1223 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1224 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1225 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1226 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1227 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1228 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1229 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1230 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1231 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1232 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1233 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1234 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1235 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1236 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1237 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1238 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1239 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1240 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1241 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1242 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1243 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1244 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1245 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1246 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1247 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1248 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1249 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1250 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1251 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1252 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1253 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1254 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1255 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1256 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1257 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1258 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1259 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1260 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1261 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1262 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1263 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1264 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1265 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1266 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1267 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1268 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1269 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1270 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1271 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1272 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1273 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1274 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1275 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1276 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1277 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1278 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1279 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1280 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1281 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1282 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1283 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1284 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1285 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1286 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1287 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1288 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1289 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1290 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1291 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1292 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1293 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1294 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1295 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1296 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1297 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1298 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1299 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1300 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1301 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1302 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1303 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1304 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1305 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1306 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1307 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1308 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1309 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1310 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1311 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1312 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1313 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1314 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1315 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1316 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1317 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1318 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1319 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1320 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1321 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1322 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1323 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1324 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1325 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1326 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1327 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1328 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1329 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1330 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1331 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1332 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1333 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1334 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1335 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1336 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1337 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1338 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1339 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1340 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1341 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1342 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1343 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1344 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1345 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1346 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1347 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1348 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1349 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1350 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1351 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1352 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1353 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1354 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1355 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1356 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1357 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1358 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1359 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1360 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1361 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1362 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1363 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1364 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1365 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1366 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1367 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1368 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1369 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1370 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1371 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1372 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1373 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1374 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1375 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1376 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1377 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1378 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1379 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1380 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1381 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1382 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1383 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1384 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1385 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1386 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1387 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1388 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1389 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1390 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1391 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1392 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1393 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1394 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1395 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1396 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1397 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1398 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1399 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1400 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1401 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1402 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1403 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1404 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1405 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1406 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1407 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1408 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1409 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1410 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1411 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1412 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1413 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1414 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1415 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1416 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1417 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1418 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1419 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1420 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1421 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1422 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1423 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1424 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1425 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1426 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1427 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1428 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1429 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1430 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1431 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1432 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1433 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1434 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1435 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1436 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1437 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1438 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1439 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1440 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1441 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1442 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1443 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1444 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1445 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1446 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1447 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1448 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1449 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1450 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1451 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1452 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1453 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1454 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1455 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1456 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1457 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1458 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1459 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1460 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1461 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1462 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1463 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1464 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1465 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1466 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1467 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1468 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1469 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1470 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1471 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1472 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1473 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1474 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1475 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1476 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1477 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1478 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1479 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1480 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1481 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1482 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1483 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1484 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1485 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1486 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1487 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1488 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1489 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1490 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1491 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1492 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1493 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1494 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1495 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1496 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1497 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1498 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1499 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1500 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1501 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1502 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1503 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1504 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1505 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1506 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1507 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1508 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1509 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1510 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1511 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1512 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1513 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1514 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1515 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1516 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1517 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1518 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1519 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1520 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1521 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1522 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1523 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1524 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1525 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1526 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1527 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1528 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1529 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1530 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1531 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1532 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1533 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1534 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1535 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1536 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1537 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1538 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1539 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1540 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1541 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1542 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1543 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1544 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1545 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1546 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1547 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1548 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1549 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1550 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1551 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1552 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1553 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1554 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1555 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1556 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1557 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1558 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1559 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1560 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1561 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1562 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1563 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1564 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1565 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1566 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1567 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1568 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1569 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1570 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1571 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1572 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1573 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1574 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1575 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1576 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1577 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1578 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1579 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1580 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1581 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1582 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1583 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1584 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1585 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1586 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1587 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1588 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1589 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1590 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1591 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1592 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1593 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1594 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1595 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1596 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1597 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1598 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1599 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1600 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1601 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1602 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1603 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1604 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1605 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1606 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1607 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1608 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1609 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1610 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1611 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1612 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1613 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1614 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1615 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1616 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1617 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1618 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1619 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1620 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1621 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1622 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1623 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1624 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1625 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1626 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1627 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1628 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1629 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1630 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1631 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1632 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1633 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1634 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1635 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1636 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1637 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1638 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1639 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1640 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1641 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1642 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1643 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1644 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1645 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1646 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1647 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1648 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1649 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1650 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1651 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1652 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1653 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1654 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1655 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1656 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1657 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1658 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1659 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1660 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1661 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1662 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1663 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1664 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1665 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1666 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1667 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1668 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1669 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1670 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1671 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1672 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1673 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1674 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1675 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1676 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1677 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1678 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1679 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1680 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1681 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1682 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1683 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1684 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1685 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1686 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1687 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1688 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1689 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1690 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1691 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1692 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1693 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1694 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1695 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1696 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1697 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1698 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1699 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1700 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1701 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1702 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1703 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1704 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1705 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1706 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1707 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1708 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1709 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1710 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1711 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1712 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1713 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1714 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1715 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1716 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1717 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1718 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1719 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1720 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1721 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1722 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1723 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1724 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1725 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1726 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1727 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1728 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1729 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1730 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1731 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1732 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1733 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1734 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1735 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1736 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1737 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1738 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1739 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1740 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1741 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1742 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1743 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1744 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1745 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1746 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1747 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1748 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1749 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1750 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1751 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1752 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1753 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1754 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1755 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1756 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1757 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1758 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1759 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1760 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1761 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1762 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1763 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1764 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1765 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1766 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1767 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1768 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1769 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1770 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1771 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1772 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1773 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1774 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1775 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1776 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1777 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1778 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1779 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1780 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1781 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1782 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1783 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1784 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1785 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1786 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1787 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1788 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1789 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1790 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1791 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1792 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1793 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1794 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1795 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1796 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1797 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1798 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1799 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1800 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1801 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1802 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1803 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1804 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1805 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1806 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1807 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1808 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1809 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1810 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1811 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1812 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1813 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1814 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1815 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1816 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1817 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1818 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1819 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1820 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1821 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1822 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1823 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1824 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1825 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1826 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1827 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1828 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1829 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1830 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1831 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1832 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1833 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1834 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1835 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1836 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1837 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1838 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1839 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1840 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1841 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1842 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1843 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1844 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1845 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1846 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1847 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1848 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1849 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1850 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1851 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1852 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1853 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1854 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1855 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1856 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1857 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1858 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1859 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1860 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1861 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1862 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1863 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1864 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1865 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1866 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1867 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1868 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1869 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1870 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1871 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1872 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1873 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1874 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1875 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1876 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1877 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1878 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1879 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1880 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1881 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1882 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1883 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1884 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1885 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1886 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1887 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1888 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1889 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1890 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1891 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1892 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1893 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1894 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1895 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1896 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1897 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1898 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1899 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1900 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1901 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1902 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		others => x"00000000"
	);


begin

	process(i_clk)
	begin
		if rising_edge(i_clk) then
			-- memory write --
			if i_we = '1' then
				mem(to_integer(unsigned(i_w_addr))) <= i_data;
			end if;
			-- memory read -- 
			o_data <= mem(to_integer(unsigned(i_r_addr)));
			
		end if; 
	end process;

end architecture arch;

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity ram is
	generic
	(
		DATA_WIDTH : natural := 32;		    -- 4 byte one line of memory
		ADDR_WIDTH : natural := 13			    -- 24576 bytes size of memory
	);

	port(
		i_clk    : in  std_logic;
		i_r_addr : in  std_logic_vector(ADDR_WIDTH-1 downto 0);
		i_data   : in  std_logic_vector(DATA_WIDTH-1 downto 0);
		i_we     : in  std_logic;
		i_w_addr : in  std_logic_vector(ADDR_WIDTH-1 downto 0);
		o_data   : out std_logic_vector(DATA_WIDTH-1 downto 0)
	);
end entity ram;

architecture arch of ram is

	type ram_t is array (0 to 2**ADDR_WIDTH-1) of std_logic_vector(DATA_WIDTH-1 downto 0);


-- GENERATED BY BC_MEM_PACKER

-- DATE: Thu May 18 16:01:02 2017

	signal mem : ram_t := (

--			***** COLOR PALLETE *****


		0 =>	x"00000000", -- R: 0 G: 0 B: 0
		1 =>	x"00C0A000", -- R: 0 G: 160 B: 192
		2 =>	x"00C0C0C0", -- R: 192 G: 192 B: 192
		3 =>	x"00C0DCC0", -- R: 192 G: 220 B: 192
		4 =>	x"00404040", -- R: 64 G: 64 B: 64
		5 =>	x"00808080", -- R: 128 G: 128 B: 128
		6 =>	x"0080A0A0", -- R: 160 G: 160 B: 128
		7 =>	x"00406080", -- R: 128 G: 96 B: 64
		8 =>	x"008080A0", -- R: 160 G: 128 B: 128
		9 =>	x"008080C0", -- R: 192 G: 128 B: 128
		10 =>	x"004060A0", -- R: 160 G: 96 B: 64
		11 =>	x"0080A0E0", -- R: 224 G: 160 B: 128
		12 =>	x"0080A0C0", -- R: 192 G: 160 B: 128
		13 =>	x"008080E0", -- R: 224 G: 128 B: 128
		14 =>	x"008060C0", -- R: 192 G: 96 B: 128
		15 =>	x"008060E0", -- R: 224 G: 96 B: 128
		16 =>	x"0080C0E0", -- R: 224 G: 192 B: 128
		17 =>	x"00A4A0A0", -- R: 160 G: 160 B: 164
		18 =>	x"00808060", -- R: 96 G: 128 B: 128
		19 =>	x"00806060", -- R: 96 G: 96 B: 128
		20 =>	x"0080A080", -- R: 128 G: 160 B: 128
		21 =>	x"00C0A080", -- R: 128 G: 160 B: 192
		22 =>	x"00C0A060", -- R: 96 G: 160 B: 192
		23 =>	x"00806040", -- R: 64 G: 96 B: 128
		24 =>	x"00806020", -- R: 32 G: 96 B: 128
		25 =>	x"00406060", -- R: 96 G: 96 B: 64
		26 =>	x"00004080", -- R: 128 G: 64 B: 0
		27 =>	x"00404060", -- R: 96 G: 64 B: 64
		28 =>	x"00006080", -- R: 128 G: 96 B: 0
		29 =>	x"00004060", -- R: 96 G: 64 B: 0
		30 =>	x"00002040", -- R: 64 G: 32 B: 0
		31 =>	x"00404080", -- R: 128 G: 64 B: 64
		32 =>	x"004060C0", -- R: 192 G: 96 B: 64
		33 =>	x"00FEFCFA", -- R: 250 G: 252 B: 254
		34 =>	x"00FDFAF7", -- R: 247 G: 250 B: 253
		35 =>	x"00FDFBF9", -- R: 249 G: 251 B: 253
		36 =>	x"00FEFDFC", -- R: 252 G: 253 B: 254
		37 =>	x"00FBF9F7", -- R: 247 G: 249 B: 251
		38 =>	x"00FDF8F5", -- R: 245 G: 248 B: 253
		39 =>	x"00FEFEFE", -- R: 254 G: 254 B: 254
		40 =>	x"00FCF6F2", -- R: 242 G: 246 B: 252
		41 =>	x"00FDFCFA", -- R: 250 G: 252 B: 253
		42 =>	x"00FEFDFB", -- R: 251 G: 253 B: 254
		43 =>	x"00FFFFFE", -- R: 254 G: 255 B: 255
		44 =>	x"00E8E0D7", -- R: 215 G: 224 B: 232
		45 =>	x"00DAD1C5", -- R: 197 G: 209 B: 218
		46 =>	x"00E6DBD0", -- R: 208 G: 219 B: 230
		47 =>	x"00FAEEE6", -- R: 230 G: 238 B: 250
		48 =>	x"00FAF6F2", -- R: 242 G: 246 B: 250
		49 =>	x"00FBF1EA", -- R: 234 G: 241 B: 251
		50 =>	x"00FFFEFD", -- R: 253 G: 254 B: 255
		51 =>	x"00FFFFFF", -- R: 255 G: 255 B: 255
		52 =>	x"00FCFBF9", -- R: 249 G: 251 B: 252
		53 =>	x"00FBF7F3", -- R: 243 G: 247 B: 251
		54 =>	x"00D9D3C8", -- R: 200 G: 211 B: 217
		55 =>	x"00CAC2B3", -- R: 179 G: 194 B: 202
		56 =>	x"00E0D6CB", -- R: 203 G: 214 B: 224
		57 =>	x"00F3E7DF", -- R: 223 G: 231 B: 243
		58 =>	x"00EFE6DE", -- R: 222 G: 230 B: 239
		59 =>	x"00F2EBE5", -- R: 229 G: 235 B: 242
		60 =>	x"00F0E5DC", -- R: 220 G: 229 B: 240
		61 =>	x"00FDFBF8", -- R: 248 G: 251 B: 253
		62 =>	x"00FFFFFD", -- R: 253 G: 255 B: 255
		63 =>	x"00FAF3ED", -- R: 237 G: 243 B: 250
		64 =>	x"00FDF9F7", -- R: 247 G: 249 B: 253
		65 =>	x"00F0EBE5", -- R: 229 G: 235 B: 240
		66 =>	x"00CBC4B7", -- R: 183 G: 196 B: 203
		67 =>	x"00D1C9BB", -- R: 187 G: 201 B: 209
		68 =>	x"00E8DDD3", -- R: 211 G: 221 B: 232
		69 =>	x"00EDE1D8", -- R: 216 G: 225 B: 237
		70 =>	x"00E6DBD1", -- R: 209 G: 219 B: 230
		71 =>	x"00DDD3C7", -- R: 199 G: 211 B: 221
		72 =>	x"00DAD0C3", -- R: 195 G: 208 B: 218
		73 =>	x"00FBF4EF", -- R: 239 G: 244 B: 251
		74 =>	x"00FFFDF9", -- R: 249 G: 253 B: 255
		75 =>	x"00FFFDFB", -- R: 251 G: 253 B: 255
		76 =>	x"00FEF7F2", -- R: 242 G: 247 B: 254
		77 =>	x"00F7ECE6", -- R: 230 G: 236 B: 247
		78 =>	x"00F6EFEB", -- R: 235 G: 239 B: 246
		79 =>	x"00E1DAD0", -- R: 208 G: 218 B: 225
		80 =>	x"00C9C0B2", -- R: 178 G: 192 B: 201
		81 =>	x"00D9D0C4", -- R: 196 G: 208 B: 217
		82 =>	x"00DED4C8", -- R: 200 G: 212 B: 222
		83 =>	x"00E4DACF", -- R: 207 G: 218 B: 228
		84 =>	x"00DFD5CA", -- R: 202 G: 213 B: 223
		85 =>	x"00DCD1C6", -- R: 198 G: 209 B: 220
		86 =>	x"00F7ECE4", -- R: 228 G: 236 B: 247
		87 =>	x"00FDF2EC", -- R: 236 G: 242 B: 253
		88 =>	x"00FDF4EE", -- R: 238 G: 244 B: 253
		89 =>	x"00FFFCF8", -- R: 248 G: 252 B: 255
		90 =>	x"00FEF6F1", -- R: 241 G: 246 B: 254
		91 =>	x"00FBF0E9", -- R: 233 G: 240 B: 251
		92 =>	x"00F9F0EB", -- R: 235 G: 240 B: 249
		93 =>	x"00F1EEEA", -- R: 234 G: 238 B: 241
		94 =>	x"00CEC5B7", -- R: 183 G: 197 B: 206
		95 =>	x"00E1D7CC", -- R: 204 G: 215 B: 225
		96 =>	x"00E7DCD1", -- R: 209 G: 220 B: 231
		97 =>	x"00ECE1D8", -- R: 216 G: 225 B: 236
		98 =>	x"00EBE0D7", -- R: 215 G: 224 B: 235
		99 =>	x"00CFC7B9", -- R: 185 G: 199 B: 207
		100 =>	x"00DCD2C7", -- R: 199 G: 210 B: 220
		101 =>	x"00F1E4DC", -- R: 220 G: 228 B: 241
		102 =>	x"00FEF2EC", -- R: 236 G: 242 B: 254
		103 =>	x"00FCF1EB", -- R: 235 G: 241 B: 252
		104 =>	x"00F6EAE3", -- R: 227 G: 234 B: 246
		105 =>	x"00F5EAE3", -- R: 227 G: 234 B: 245
		106 =>	x"00FDFBFA", -- R: 250 G: 251 B: 253
		107 =>	x"00D9D0C5", -- R: 197 G: 208 B: 217
		108 =>	x"00DFD5C9", -- R: 201 G: 213 B: 223
		109 =>	x"00F2E7DE", -- R: 222 G: 231 B: 242
		110 =>	x"00ECE0D7", -- R: 215 G: 224 B: 236
		111 =>	x"00E2D8CD", -- R: 205 G: 216 B: 226
		112 =>	x"00D6CDC1", -- R: 193 G: 205 B: 214
		113 =>	x"00BFB9A9", -- R: 169 G: 185 B: 191
		114 =>	x"00C7C0B1", -- R: 177 G: 192 B: 199
		115 =>	x"00CCC4B6", -- R: 182 G: 196 B: 204
		116 =>	x"00EDE1D9", -- R: 217 G: 225 B: 237
		117 =>	x"00F9ECE6", -- R: 230 G: 236 B: 249
		118 =>	x"00F6EAE2", -- R: 226 G: 234 B: 246
		119 =>	x"00E9DED5", -- R: 213 G: 222 B: 233
		120 =>	x"00F8F4F1", -- R: 241 G: 244 B: 248
		121 =>	x"00FAF8F7", -- R: 247 G: 248 B: 250
		122 =>	x"00DCD3C7", -- R: 199 G: 211 B: 220
		123 =>	x"00E3D9CE", -- R: 206 G: 217 B: 227
		124 =>	x"00C7C1B1", -- R: 177 G: 193 B: 199
		125 =>	x"00B8B3A3", -- R: 163 G: 179 B: 184
		126 =>	x"00B0AC9B", -- R: 155 G: 172 B: 176
		127 =>	x"00B4AF9E", -- R: 158 G: 175 B: 180
		128 =>	x"00B9B3A3", -- R: 163 G: 179 B: 185
		129 =>	x"00C4BDAE", -- R: 174 G: 189 B: 196
		130 =>	x"00F1E5DD", -- R: 221 G: 229 B: 241
		131 =>	x"00F3E8E0", -- R: 224 G: 232 B: 243
		132 =>	x"00DFD4C9", -- R: 201 G: 212 B: 223
		133 =>	x"00EBE4DD", -- R: 221 G: 228 B: 235
		134 =>	x"00E2DCD4", -- R: 212 G: 220 B: 226
		135 =>	x"00D3C9BB", -- R: 187 G: 201 B: 211
		136 =>	x"00CCC3B5", -- R: 181 G: 195 B: 204
		137 =>	x"00B6B1A0", -- R: 160 G: 177 B: 182
		138 =>	x"00AEAA99", -- R: 153 G: 170 B: 174
		139 =>	x"00ABA796", -- R: 150 G: 167 B: 171
		140 =>	x"00B0AC9A", -- R: 154 G: 172 B: 176
		141 =>	x"00B5B09F", -- R: 159 G: 176 B: 181
		142 =>	x"00BBB6A6", -- R: 166 G: 182 B: 187
		143 =>	x"00C7BFB1", -- R: 177 G: 191 B: 199
		144 =>	x"00D6CCC0", -- R: 192 G: 204 B: 214
		145 =>	x"00E1D7CB", -- R: 203 G: 215 B: 225
		146 =>	x"00D7CEC1", -- R: 193 G: 206 B: 215
		147 =>	x"00EEEAE4", -- R: 228 G: 234 B: 238
		148 =>	x"00F3EFEB", -- R: 235 G: 239 B: 243
		149 =>	x"00E1D9CF", -- R: 207 G: 217 B: 225
		150 =>	x"00C2BDAD", -- R: 173 G: 189 B: 194
		151 =>	x"00B1AC9B", -- R: 155 G: 172 B: 177
		152 =>	x"00AFAB99", -- R: 153 G: 171 B: 175
		153 =>	x"00B2AE9C", -- R: 156 G: 174 B: 178
		154 =>	x"00BDB7A7", -- R: 167 G: 183 B: 189
		155 =>	x"00CAC2B4", -- R: 180 G: 194 B: 202
		156 =>	x"00DAD1C4", -- R: 196 G: 209 B: 218
		157 =>	x"00EBE7E1", -- R: 225 G: 231 B: 235
		158 =>	x"00BEB8A8", -- R: 168 G: 184 B: 190
		159 =>	x"00B0AB9A", -- R: 154 G: 171 B: 176
		160 =>	x"00A5A290", -- R: 144 G: 162 B: 165
		161 =>	x"00ADA998", -- R: 152 G: 169 B: 173
		162 =>	x"00BBB5A5", -- R: 165 G: 181 B: 187
		163 =>	x"00C8C0B2", -- R: 178 G: 192 B: 200
		164 =>	x"00DCD3C8", -- R: 200 G: 211 B: 220
		165 =>	x"00E3D8CE", -- R: 206 G: 216 B: 227
		166 =>	x"00E2DACF", -- R: 207 G: 218 B: 226
		167 =>	x"00DCD5CA", -- R: 202 G: 213 B: 220
		168 =>	x"00B9B2A0", -- R: 160 G: 178 B: 185
		169 =>	x"00BCB5A5", -- R: 165 G: 181 B: 188
		170 =>	x"00B6B19F", -- R: 159 G: 177 B: 182
		171 =>	x"00BAB3A2", -- R: 162 G: 179 B: 186
		172 =>	x"00BFB8A9", -- R: 169 G: 184 B: 191
		173 =>	x"00DBD2C6", -- R: 198 G: 210 B: 219
		174 =>	x"00EFE9E4", -- R: 228 G: 233 B: 239
		175 =>	x"00ECE8E2", -- R: 226 G: 232 B: 236
		176 =>	x"00F1EDE8", -- R: 232 G: 237 B: 241
		177 =>	x"00EFEBE6", -- R: 230 G: 235 B: 239
		178 =>	x"00DBD5CC", -- R: 204 G: 213 B: 219
		179 =>	x"00C9C1B2", -- R: 178 G: 193 B: 201
		180 =>	x"00CBC3B5", -- R: 181 G: 195 B: 203
		181 =>	x"00DDD6CC", -- R: 204 G: 214 B: 221
		182 =>	x"00E4DDD4", -- R: 212 G: 221 B: 228
		183 =>	x"00F9F6F4", -- R: 244 G: 246 B: 249
		184 =>	x"00F6F3EF", -- R: 239 G: 243 B: 246
		185 =>	x"00FFFEFE", -- R: 254 G: 254 B: 255
		186 =>	x"004CB122", -- R: 34 G: 177 B: 76
		187 =>	x"003D8B1B", -- R: 27 G: 139 B: 61
		188 =>	x"001DE6B5", -- R: 181 G: 230 B: 29
		189 =>	x"008060A0", -- R: 160 G: 96 B: 128
		190 =>	x"00002060", -- R: 96 G: 32 B: 0
		191 =>	x"00402060", -- R: 96 G: 32 B: 64
		192 =>	x"00888888", -- R: 136 G: 136 B: 136
		193 =>	x"00777777", -- R: 119 G: 119 B: 119
		194 =>	x"00999999", -- R: 153 G: 153 B: 153
		195 =>	x"00666666", -- R: 102 G: 102 B: 102
		196 =>	x"00AAAAAA", -- R: 170 G: 170 B: 170
		197 =>	x"00555555", -- R: 85 G: 85 B: 85
		198 =>	x"00BBBBBB", -- R: 187 G: 187 B: 187
		199 =>	x"00444444", -- R: 68 G: 68 B: 68
		200 =>	x"00333333", -- R: 51 G: 51 B: 51
		201 =>	x"00222222", -- R: 34 G: 34 B: 34
		202 =>	x"00111111", -- R: 17 G: 17 B: 17
		203 =>	x"00CCCCCC", -- R: 204 G: 204 B: 204
		204 =>	x"004080A0", -- R: 160 G: 128 B: 64
		205 =>	x"00000000", -- Unused
		206 =>	x"00000000", -- Unused
		207 =>	x"00000000", -- Unused
		208 =>	x"00000000", -- Unused
		209 =>	x"00000000", -- Unused
		210 =>	x"00000000", -- Unused
		211 =>	x"00000000", -- Unused
		212 =>	x"00000000", -- Unused
		213 =>	x"00000000", -- Unused
		214 =>	x"00000000", -- Unused
		215 =>	x"00000000", -- Unused
		216 =>	x"00000000", -- Unused
		217 =>	x"00000000", -- Unused
		218 =>	x"00000000", -- Unused
		219 =>	x"00000000", -- Unused
		220 =>	x"00000000", -- Unused
		221 =>	x"00000000", -- Unused
		222 =>	x"00000000", -- Unused
		223 =>	x"00000000", -- Unused
		224 =>	x"00000000", -- Unused
		225 =>	x"00000000", -- Unused
		226 =>	x"00000000", -- Unused
		227 =>	x"00000000", -- Unused
		228 =>	x"00000000", -- Unused
		229 =>	x"00000000", -- Unused
		230 =>	x"00000000", -- Unused
		231 =>	x"00000000", -- Unused
		232 =>	x"00000000", -- Unused
		233 =>	x"00000000", -- Unused
		234 =>	x"00000000", -- Unused
		235 =>	x"00000000", -- Unused
		236 =>	x"00000000", -- Unused
		237 =>	x"00000000", -- Unused
		238 =>	x"00000000", -- Unused
		239 =>	x"00000000", -- Unused
		240 =>	x"00000000", -- Unused
		241 =>	x"00000000", -- Unused
		242 =>	x"00000000", -- Unused
		243 =>	x"00000000", -- Unused
		244 =>	x"00000000", -- Unused
		245 =>	x"00000000", -- Unused
		246 =>	x"00000000", -- Unused
		247 =>	x"00000000", -- Unused
		248 =>	x"00000000", -- Unused
		249 =>	x"00000000", -- Unused
		250 =>	x"00000000", -- Unused
		251 =>	x"00000000", -- Unused
		252 =>	x"00000000", -- Unused
		253 =>	x"00000000", -- Unused
		254 =>	x"00000000", -- Unused

--			***** 16x16 IMAGES *****




		255 =>	x"01010101", -- IMG_16x18_crvcina_desno
		256 =>	x"01010101",
		257 =>	x"01020101",
		258 =>	x"01010101",
		259 =>	x"01010101",
		260 =>	x"01010301",
		261 =>	x"04040101",
		262 =>	x"01010101",
		263 =>	x"01010101",
		264 =>	x"01050006",
		265 =>	x"07080101",
		266 =>	x"01010101",
		267 =>	x"01010101",
		268 =>	x"02090A0B",
		269 =>	x"0B0C0101",
		270 =>	x"01010101",
		271 =>	x"0101010C",
		272 =>	x"0D0B0B0B",
		273 =>	x"0B0B0201",
		274 =>	x"01010101",
		275 =>	x"0101010E",
		276 =>	x"0D0D0B0B",
		277 =>	x"0D0B0201",
		278 =>	x"01010101",
		279 =>	x"01010109",
		280 =>	x"0F0D0202",
		281 =>	x"0B020201",
		282 =>	x"03050101",
		283 =>	x"01010102",
		284 =>	x"0E0D0B10",
		285 =>	x"0B0B1103",
		286 =>	x"05121314",
		287 =>	x"01010101",
		288 =>	x"0C0E0811",
		289 =>	x"11111115",
		290 =>	x"16121705",
		291 =>	x"01010202",
		292 =>	x"02051812",
		293 =>	x"12191A1B",
		294 =>	x"12121101",
		295 =>	x"01071A1C",
		296 =>	x"1A121515",
		297 =>	x"171D1A07",
		298 =>	x"19110101",
		299 =>	x"01071A1D",
		300 =>	x"1E1F0908",
		301 =>	x"1B200E09",
		302 =>	x"02010101",
		303 =>	x"01191E1E",
		304 =>	x"1F0F0F0D",
		305 =>	x"0B0D0902",
		306 =>	x"01010101",
		307 =>	x"11191E07",
		308 =>	x"0E0E0A09",
		309 =>	x"0B0C0C01",
		310 =>	x"01010101",
		311 =>	x"01020202",
		312 =>	x"02020202",
		313 =>	x"02020201",
		314 =>	x"01010101",
		315 =>	x"01030202",
		316 =>	x"03030203",
		317 =>	x"02030301",
		318 =>	x"01010101",
		319 =>	x"01010101", -- IMG_16x18_crvcina_levo
		320 =>	x"01010201",
		321 =>	x"01010101",
		322 =>	x"01010101",
		323 =>	x"01010101",
		324 =>	x"01010404",
		325 =>	x"01030101",
		326 =>	x"01010101",
		327 =>	x"01010101",
		328 =>	x"01010807",
		329 =>	x"06000501",
		330 =>	x"01010101",
		331 =>	x"01010101",
		332 =>	x"01010C0B",
		333 =>	x"0B0A0902",
		334 =>	x"01010101",
		335 =>	x"01010101",
		336 =>	x"01020B0B",
		337 =>	x"0B0B0B0D",
		338 =>	x"0C010101",
		339 =>	x"01010101",
		340 =>	x"01020B0D",
		341 =>	x"0B0B0D0D",
		342 =>	x"0E010101",
		343 =>	x"01010503",
		344 =>	x"0102020B",
		345 =>	x"02020D0F",
		346 =>	x"09010101",
		347 =>	x"14131205",
		348 =>	x"03110B0B",
		349 =>	x"100B0D0E",
		350 =>	x"02010101",
		351 =>	x"05171216",
		352 =>	x"15111111",
		353 =>	x"11080E0C",
		354 =>	x"01010101",
		355 =>	x"01111212",
		356 =>	x"1B1A1912",
		357 =>	x"12180502",
		358 =>	x"02020101",
		359 =>	x"01011119",
		360 =>	x"071A1D17",
		361 =>	x"1515121A",
		362 =>	x"1C1A0701",
		363 =>	x"01010102",
		364 =>	x"090E201B",
		365 =>	x"08091F1E",
		366 =>	x"1D1A0701",
		367 =>	x"01010101",
		368 =>	x"02090D0B",
		369 =>	x"0D0F0F1F",
		370 =>	x"1E1E1901",
		371 =>	x"01010101",
		372 =>	x"020C0C0B",
		373 =>	x"090A0E0E",
		374 =>	x"071E1911",
		375 =>	x"01010101",
		376 =>	x"01020202",
		377 =>	x"02020202",
		378 =>	x"02020201",
		379 =>	x"01010101",
		380 =>	x"01030302",
		381 =>	x"03020303",
		382 =>	x"02020301",
		383 =>	x"01010101", -- IMG_16x18_nebo_svetlo
		384 =>	x"01010101",
		385 =>	x"01010101",
		386 =>	x"01010101",
		387 =>	x"01010101",
		388 =>	x"01010101",
		389 =>	x"01010101",
		390 =>	x"01010101",
		391 =>	x"01010101",
		392 =>	x"01010101",
		393 =>	x"01010101",
		394 =>	x"01010101",
		395 =>	x"01010101",
		396 =>	x"01010101",
		397 =>	x"01010101",
		398 =>	x"01010101",
		399 =>	x"01010101",
		400 =>	x"01010101",
		401 =>	x"01010101",
		402 =>	x"01010101",
		403 =>	x"01010101",
		404 =>	x"01010101",
		405 =>	x"01010101",
		406 =>	x"01010101",
		407 =>	x"01010101",
		408 =>	x"01010101",
		409 =>	x"01010101",
		410 =>	x"01010101",
		411 =>	x"01010101",
		412 =>	x"01010101",
		413 =>	x"01010101",
		414 =>	x"01010101",
		415 =>	x"01010101",
		416 =>	x"01010101",
		417 =>	x"01010101",
		418 =>	x"01010101",
		419 =>	x"01010101",
		420 =>	x"01010101",
		421 =>	x"01010101",
		422 =>	x"01010101",
		423 =>	x"01010101",
		424 =>	x"01010101",
		425 =>	x"01010101",
		426 =>	x"01010101",
		427 =>	x"01010101",
		428 =>	x"01010101",
		429 =>	x"01010101",
		430 =>	x"01010101",
		431 =>	x"01010101",
		432 =>	x"01010101",
		433 =>	x"01010101",
		434 =>	x"01010101",
		435 =>	x"01010101",
		436 =>	x"01010101",
		437 =>	x"01010101",
		438 =>	x"01010101",
		439 =>	x"01010101",
		440 =>	x"01010101",
		441 =>	x"01010101",
		442 =>	x"01010101",
		443 =>	x"01010101",
		444 =>	x"01010101",
		445 =>	x"01010101",
		446 =>	x"01010101",
		447 =>	x"01010101", -- IMG_16x18_oblak
		448 =>	x"01010101",
		449 =>	x"01010101",
		450 =>	x"01010101",
		451 =>	x"01010101",
		452 =>	x"01010121",
		453 =>	x"22230101",
		454 =>	x"01010101",
		455 =>	x"01242526",
		456 =>	x"01012728",
		457 =>	x"292A2A01",
		458 =>	x"01010101",
		459 =>	x"2B2C2D2E",
		460 =>	x"2F013031",
		461 =>	x"2B323334",
		462 =>	x"35010101",
		463 =>	x"33363738",
		464 =>	x"393A3B3C",
		465 =>	x"3D3E2B24",
		466 =>	x"3F400101",
		467 =>	x"41424344",
		468 =>	x"45464748",
		469 =>	x"494A4B33",
		470 =>	x"4C4D4E01",
		471 =>	x"4F505152",
		472 =>	x"46535455",
		473 =>	x"56575859",
		474 =>	x"5A5B5C01",
		475 =>	x"5D5E5F46",
		476 =>	x"60616263",
		477 =>	x"64606566",
		478 =>	x"67686901",
		479 =>	x"6A6B6C6D",
		480 =>	x"6E6F7071",
		481 =>	x"72732D74",
		482 =>	x"75767778",
		483 =>	x"33797A7B",
		484 =>	x"7A7C7D7E",
		485 =>	x"7F808170",
		486 =>	x"82838485",
		487 =>	x"01018687",
		488 =>	x"88898A8B",
		489 =>	x"8C8D8E8F",
		490 =>	x"90919293",
		491 =>	x"01019495",
		492 =>	x"3696978B",
		493 =>	x"98999A9B",
		494 =>	x"9C2E5F01",
		495 =>	x"01010101",
		496 =>	x"9D9E9FA0",
		497 =>	x"A199A2A3",
		498 =>	x"A4A5A632",
		499 =>	x"01010101",
		500 =>	x"A7A8A9AA",
		501 =>	x"AB9A9EAC",
		502 =>	x"50ADAE01",
		503 =>	x"01010101",
		504 =>	x"01AFB0B1",
		505 =>	x"B2B3B4B5",
		506 =>	x"B6B70101",
		507 =>	x"01010101",
		508 =>	x"01010101",
		509 =>	x"01B8B8B9",
		510 =>	x"01010101",
		511 =>	x"BABABBBA", -- IMG_16x18_tobla1
		512 =>	x"BABABABA",
		513 =>	x"BBBABABB",
		514 =>	x"BBBBBBBB",
		515 =>	x"BBBBBBBB",
		516 =>	x"BBBBBABA",
		517 =>	x"BCBBBBBA",
		518 =>	x"BBBABBBA",
		519 =>	x"BBBBBABB",
		520 =>	x"BBBABABC",
		521 =>	x"BCBCBBBA",
		522 =>	x"BBBBBBBB",
		523 =>	x"BBBBBBBB",
		524 =>	x"BBBABCBC",
		525 =>	x"BBBBBBBB",
		526 =>	x"BBBBBCBA",
		527 =>	x"BABCBBBB",
		528 =>	x"BBBBBBBB",
		529 =>	x"BCBCBBBB",
		530 =>	x"BBBCBCBC",
		531 =>	x"BCBCBCBB",
		532 =>	x"BABABBBB",
		533 =>	x"BBBBBBBB",
		534 =>	x"BBBBBCBB",
		535 =>	x"BCBABCBC",
		536 =>	x"BBBBBBBB",
		537 =>	x"BBBBBBBB",
		538 =>	x"BBBCBBBC",
		539 =>	x"BCBCBCBB",
		540 =>	x"BBBBBBBB",
		541 =>	x"BBBABBBB",
		542 =>	x"BABBBCBB",
		543 =>	x"BABCBBBB",
		544 =>	x"BBBBBABB",
		545 =>	x"BBBB0ABB",
		546 =>	x"BBBBBBBA",
		547 =>	x"BBBBBABB",
		548 =>	x"BBBCBBBB",
		549 =>	x"09BBBCBA",
		550 =>	x"BBBABB0A",
		551 =>	x"0ABABA0A",
		552 =>	x"BCBCBCBB",
		553 =>	x"BBBBBCBC",
		554 =>	x"BBBB0A0A",
		555 =>	x"BBBDBABA",
		556 =>	x"BBBCBCBB",
		557 =>	x"BABCBCBC",
		558 =>	x"BC091F1F",
		559 =>	x"BBBBBBBB",
		560 =>	x"BCBCBCBA",
		561 =>	x"BBBCBCBC",
		562 =>	x"BA091F07",
		563 =>	x"1FBBBBBB",
		564 =>	x"BBBCBABB",
		565 =>	x"0ABBBC0A",
		566 =>	x"0A090A0A",
		567 =>	x"1F0ABABA",
		568 =>	x"BABABBBB",
		569 =>	x"BBBEBB0A",
		570 =>	x"0A0A0ABF",
		571 =>	x"0A09BD1F",
		572 =>	x"BA090A0A",
		573 =>	x"BB0A090A",
		574 =>	x"0A0A0707",
		575 =>	x"C0C1C2C2", -- IMG_16x18_tobla2
		576 =>	x"C1C1C0C0",
		577 =>	x"C3C3C0C4",
		578 =>	x"C2C0C2C1",
		579 =>	x"C1C0C3C5",
		580 =>	x"C6C0C0C1",
		581 =>	x"C1C3C7C7",
		582 =>	x"C1C7C5C5",
		583 =>	x"C5C0C1C3",
		584 =>	x"C5C3C5C0",
		585 =>	x"C0C5C3C3",
		586 =>	x"C8C5C1C0",
		587 =>	x"C7C1C2C3",
		588 =>	x"C3C1C3C5",
		589 =>	x"C0C5C7C5",
		590 =>	x"C5C8C3C7",
		591 =>	x"C3C1C3C0",
		592 =>	x"C3C3C3C7",
		593 =>	x"C5C5C3C5",
		594 =>	x"C5C1C2C0",
		595 =>	x"C8C1C1C3",
		596 =>	x"C1C5C1C5",
		597 =>	x"C1C5C2C4",
		598 =>	x"C4C4C3C0",
		599 =>	x"C1C5C3C0",
		600 =>	x"C3C3C3C3",
		601 =>	x"C1C2C1C3",
		602 =>	x"C2C3C3C0",
		603 =>	x"C7C7C1C0",
		604 =>	x"C1C9C8C5",
		605 =>	x"C8C1C3C5",
		606 =>	x"C5C3C0C1",
		607 =>	x"C3C7C9C8",
		608 =>	x"C7C5C0C1",
		609 =>	x"C8C8C5C5",
		610 =>	x"C7C1C0C7",
		611 =>	x"C2C1C7C3",
		612 =>	x"C3C1C5C1",
		613 =>	x"C5C5C1C5",
		614 =>	x"C5C0C3C5",
		615 =>	x"C3C3C9C5",
		616 =>	x"C3C7C1C4",
		617 =>	x"C0C3C9C3",
		618 =>	x"C4C0C5C3",
		619 =>	x"C5C1C5CA",
		620 =>	x"C3C5C7C5",
		621 =>	x"C9C7C5C1",
		622 =>	x"C0C3C1C1",
		623 =>	x"C0C0C2C3",
		624 =>	x"C0C1C7C7",
		625 =>	x"C5C3C8C2",
		626 =>	x"C5C2C1C7",
		627 =>	x"C2C6C2C2",
		628 =>	x"C2C5C2CB",
		629 =>	x"C2CBC2C4",
		630 =>	x"C0C0C0C7",
		631 =>	x"C3C4C6C4",
		632 =>	x"C0C5C5C5",
		633 =>	x"C1C5C4C6",
		634 =>	x"C3C8C7C1",
		635 =>	x"C2C0C4C4",
		636 =>	x"C2C800C7",
		637 =>	x"C5C9C1C3",
		638 =>	x"C7C9C3C2",
		639 =>	x"1E1B1F07", -- IMG_16x18_tobla3
		640 =>	x"070ACC0A",
		641 =>	x"0ACCCC07",
		642 =>	x"07071B1E",
		643 =>	x"1B1B0707",
		644 =>	x"CC0808CC",
		645 =>	x"0808CC07",
		646 =>	x"07071B1B",
		647 =>	x"1B070707",
		648 =>	x"CCCC08CC",
		649 =>	x"09CC0707",
		650 =>	x"0A07071B",
		651 =>	x"1B0707CC",
		652 =>	x"CC0ACCCC",
		653 =>	x"CC0808CC",
		654 =>	x"07071B1B",
		655 =>	x"1B1B07CC",
		656 =>	x"CCCCCC08",
		657 =>	x"08080A07",
		658 =>	x"CC0A1B1D",
		659 =>	x"1B0707CC",
		660 =>	x"CCCC080C",
		661 =>	x"0808CC07",
		662 =>	x"CC07071B",
		663 =>	x"1B07070A",
		664 =>	x"0ACC0809",
		665 =>	x"0C090A07",
		666 =>	x"CC071B1B",
		667 =>	x"1B07070A",
		668 =>	x"CC080908",
		669 =>	x"080808CC",
		670 =>	x"08070707",
		671 =>	x"070ACCCC",
		672 =>	x"CC080908",
		673 =>	x"080808CC",
		674 =>	x"CC07071B",
		675 =>	x"1B070ACC",
		676 =>	x"08080908",
		677 =>	x"090808CC",
		678 =>	x"080A071D",
		679 =>	x"1B070ACC",
		680 =>	x"08080808",
		681 =>	x"08CCCC08",
		682 =>	x"CC07071F",
		683 =>	x"1B0707CC",
		684 =>	x"08CC0808",
		685 =>	x"08CC07CC",
		686 =>	x"CC070707",
		687 =>	x"1D1B07CC",
		688 =>	x"CCCC0808",
		689 =>	x"CC08CC0A",
		690 =>	x"071B1B1B",
		691 =>	x"1D1B070A",
		692 =>	x"CC0808CC",
		693 =>	x"CC0A0707",
		694 =>	x"07071B1E",
		695 =>	x"1D1B1F07",
		696 =>	x"CC0808CC",
		697 =>	x"0A070707",
		698 =>	x"071B1B1D",
		699 =>	x"1E1D1B07",
		700 =>	x"0A0809CC",
		701 =>	x"CCCC071B",
		702 =>	x"071B1B1D",


--			***** MAP *****


		703 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		704 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		705 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		706 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		707 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		708 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		709 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		710 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		711 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		712 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		713 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		714 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		715 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		716 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		717 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		718 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		719 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		720 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		721 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		722 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		723 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		724 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		725 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		726 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		727 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		728 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		729 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		730 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		731 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		732 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		733 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		734 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		735 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		736 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		737 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		738 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		739 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		740 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		741 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		742 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		743 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		744 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		745 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		746 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		747 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		748 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		749 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		750 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		751 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		752 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		753 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		754 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		755 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		756 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		757 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		758 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		759 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		760 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		761 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		762 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		763 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		764 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		765 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		766 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		767 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		768 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		769 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		770 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		771 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		772 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		773 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		774 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		775 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		776 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		777 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		778 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		779 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		780 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		781 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		782 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		783 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		784 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		785 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		786 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		787 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		788 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		789 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		790 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		791 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		792 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		793 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		794 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		795 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		796 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		797 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		798 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		799 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		800 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		801 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		802 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		803 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		804 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		805 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		806 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		807 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		808 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		809 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		810 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		811 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		812 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		813 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		814 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		815 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		816 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		817 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		818 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		819 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		820 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		821 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		822 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		823 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		824 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		825 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		826 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		827 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		828 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		829 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		830 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		831 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		832 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		833 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		834 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		835 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		836 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		837 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		838 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		839 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		840 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		841 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		842 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		843 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		844 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		845 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		846 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		847 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		848 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		849 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		850 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		851 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		852 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		853 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		854 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		855 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		856 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		857 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		858 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		859 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		860 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		861 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		862 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		863 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		864 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		865 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		866 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		867 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		868 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		869 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		870 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		871 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		872 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		873 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		874 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		875 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		876 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		877 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		878 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		879 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		880 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		881 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		882 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		883 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		884 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		885 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		886 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		887 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		888 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		889 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		890 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		891 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		892 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		893 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		894 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		895 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		896 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		897 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		898 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		899 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		900 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		901 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		902 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		903 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		904 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		905 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		906 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		907 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		908 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		909 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		910 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		911 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		912 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		913 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		914 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		915 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		916 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		917 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		918 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		919 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		920 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		921 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		922 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		923 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		924 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		925 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		926 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		927 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		928 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		929 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		930 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		931 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		932 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		933 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		934 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		935 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		936 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		937 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		938 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		939 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		940 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		941 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		942 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		943 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		944 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		945 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		946 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		947 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		948 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		949 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		950 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		951 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		952 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		953 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		954 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		955 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		956 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		957 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		958 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		959 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		960 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		961 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		962 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		963 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		964 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		965 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		966 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		967 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		968 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		969 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		970 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		971 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		972 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		973 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		974 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		975 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		976 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		977 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		978 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		979 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		980 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		981 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		982 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		983 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		984 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		985 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		986 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		987 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		988 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		989 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		990 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		991 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		992 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		993 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		994 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		995 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		996 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		997 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		998 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		999 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1000 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1001 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1002 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1003 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1004 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1005 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1006 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1007 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1008 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1009 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1010 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1011 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1012 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1013 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1014 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1015 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1016 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1017 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1018 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1019 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1020 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1021 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1022 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1023 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1024 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1025 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1026 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1027 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1028 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1029 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1030 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1031 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1032 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1033 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1034 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1035 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1036 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1037 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1038 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1039 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1040 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1041 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1042 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1043 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1044 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1045 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1046 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1047 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1048 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1049 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1050 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1051 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1052 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1053 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1054 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1055 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1056 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1057 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1058 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1059 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1060 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1061 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1062 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1063 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1064 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1065 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1066 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1067 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1068 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1069 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1070 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1071 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1072 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1073 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1074 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1075 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1076 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1077 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1078 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1079 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1080 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1081 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1082 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1083 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1084 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1085 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1086 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1087 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1088 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1089 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1090 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1091 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1092 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1093 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1094 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1095 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1096 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1097 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1098 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1099 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1100 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1101 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1102 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1103 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1104 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1105 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1106 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1107 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1108 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1109 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1110 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1111 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1112 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1113 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1114 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1115 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1116 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1117 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1118 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1119 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1120 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1121 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1122 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1123 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1124 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1125 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1126 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1127 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1128 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1129 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1130 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1131 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1132 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1133 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1134 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1135 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1136 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1137 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1138 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1139 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1140 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1141 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1142 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1143 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1144 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1145 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1146 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1147 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1148 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1149 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1150 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1151 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1152 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1153 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1154 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1155 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1156 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1157 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1158 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1159 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1160 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1161 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1162 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1163 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1164 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1165 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1166 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1167 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1168 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1169 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1170 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1171 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1172 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1173 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1174 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1175 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1176 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1177 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1178 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1179 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1180 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1181 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1182 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1183 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1184 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1185 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1186 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1187 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1188 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1189 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1190 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1191 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1192 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1193 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1194 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1195 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1196 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1197 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1198 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1199 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1200 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1201 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1202 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1203 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1204 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1205 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1206 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1207 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1208 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1209 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1210 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1211 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1212 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1213 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1214 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1215 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1216 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1217 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1218 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1219 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1220 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1221 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1222 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1223 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1224 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1225 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1226 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1227 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1228 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1229 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1230 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1231 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1232 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1233 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1234 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1235 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1236 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1237 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1238 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1239 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1240 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1241 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1242 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1243 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1244 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1245 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1246 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1247 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1248 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1249 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1250 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1251 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1252 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1253 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1254 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1255 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1256 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1257 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1258 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1259 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1260 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1261 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1262 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1263 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1264 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1265 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1266 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1267 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1268 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1269 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1270 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1271 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1272 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1273 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1274 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1275 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1276 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1277 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1278 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1279 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1280 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1281 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1282 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1283 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1284 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1285 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1286 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1287 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1288 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1289 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1290 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1291 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1292 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1293 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1294 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1295 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1296 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1297 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1298 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1299 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1300 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1301 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1302 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1303 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1304 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1305 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1306 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1307 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1308 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1309 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1310 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1311 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1312 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1313 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1314 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1315 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1316 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1317 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1318 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1319 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1320 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1321 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1322 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1323 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1324 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1325 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1326 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1327 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1328 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1329 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1330 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1331 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1332 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1333 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1334 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1335 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1336 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1337 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1338 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1339 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1340 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1341 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1342 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1343 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1344 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1345 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1346 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1347 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1348 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1349 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1350 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1351 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1352 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1353 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1354 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1355 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1356 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1357 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1358 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1359 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1360 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1361 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1362 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1363 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1364 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1365 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1366 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1367 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1368 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1369 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1370 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1371 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1372 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1373 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1374 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1375 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1376 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1377 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1378 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1379 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1380 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1381 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1382 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1383 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1384 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1385 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1386 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1387 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1388 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1389 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1390 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1391 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1392 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1393 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1394 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1395 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1396 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1397 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1398 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1399 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1400 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1401 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1402 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1403 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1404 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1405 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1406 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1407 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1408 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1409 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1410 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1411 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1412 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1413 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1414 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1415 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1416 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1417 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1418 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1419 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1420 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1421 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1422 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1423 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1424 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1425 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1426 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1427 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1428 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1429 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1430 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1431 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1432 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1433 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1434 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1435 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1436 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1437 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1438 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1439 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1440 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1441 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1442 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1443 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1444 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1445 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1446 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1447 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1448 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1449 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1450 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1451 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1452 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1453 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1454 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1455 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1456 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1457 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1458 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1459 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1460 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1461 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1462 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1463 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1464 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1465 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1466 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1467 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1468 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1469 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1470 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1471 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1472 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1473 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1474 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1475 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1476 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1477 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1478 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1479 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1480 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1481 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1482 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1483 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1484 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1485 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1486 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1487 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1488 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1489 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1490 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1491 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1492 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1493 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1494 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1495 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1496 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1497 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1498 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1499 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1500 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1501 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1502 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1503 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1504 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1505 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1506 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1507 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1508 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1509 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1510 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1511 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1512 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1513 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1514 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1515 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1516 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1517 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1518 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1519 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1520 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1521 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1522 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1523 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1524 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1525 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1526 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1527 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1528 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1529 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1530 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1531 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1532 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1533 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1534 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1535 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1536 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1537 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1538 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1539 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1540 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1541 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1542 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1543 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1544 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1545 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1546 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1547 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1548 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1549 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1550 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1551 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1552 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1553 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1554 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1555 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1556 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1557 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1558 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1559 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1560 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1561 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1562 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1563 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1564 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1565 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1566 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1567 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1568 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1569 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1570 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1571 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1572 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1573 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1574 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1575 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1576 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1577 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1578 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1579 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1580 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1581 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1582 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1583 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1584 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1585 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1586 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1587 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1588 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1589 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1590 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1591 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1592 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1593 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1594 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1595 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1596 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1597 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1598 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1599 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1600 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1601 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1602 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1603 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1604 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1605 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1606 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1607 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1608 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1609 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1610 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1611 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1612 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1613 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1614 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1615 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1616 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1617 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1618 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1619 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1620 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1621 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1622 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1623 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1624 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1625 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1626 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1627 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1628 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1629 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1630 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1631 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1632 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1633 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1634 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1635 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1636 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1637 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1638 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1639 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1640 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1641 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1642 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1643 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1644 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1645 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1646 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1647 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1648 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1649 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1650 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1651 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1652 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1653 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1654 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1655 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1656 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1657 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1658 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1659 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1660 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1661 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1662 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1663 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1664 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1665 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1666 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1667 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1668 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1669 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1670 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1671 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1672 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1673 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1674 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1675 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1676 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1677 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1678 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1679 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1680 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1681 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1682 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1683 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1684 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1685 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1686 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1687 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1688 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1689 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1690 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1691 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1692 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1693 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1694 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1695 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1696 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1697 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1698 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1699 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1700 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1701 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1702 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1703 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1704 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1705 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1706 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1707 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1708 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1709 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1710 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1711 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1712 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1713 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1714 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1715 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1716 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1717 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1718 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1719 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1720 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1721 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1722 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1723 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1724 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1725 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1726 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1727 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1728 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1729 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1730 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1731 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1732 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1733 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1734 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1735 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1736 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1737 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1738 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1739 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1740 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1741 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1742 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1743 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1744 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1745 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1746 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1747 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1748 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1749 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1750 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1751 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1752 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1753 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1754 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1755 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1756 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1757 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1758 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1759 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1760 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1761 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1762 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1763 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1764 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1765 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1766 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1767 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1768 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1769 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1770 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1771 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1772 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1773 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1774 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1775 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1776 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1777 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1778 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1779 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1780 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1781 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1782 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1783 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1784 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1785 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1786 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1787 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1788 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1789 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1790 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1791 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1792 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1793 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1794 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1795 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1796 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1797 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1798 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1799 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1800 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1801 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1802 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1803 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1804 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1805 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1806 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1807 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1808 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1809 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1810 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1811 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1812 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1813 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1814 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1815 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1816 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1817 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1818 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1819 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1820 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1821 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1822 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1823 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1824 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1825 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1826 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1827 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1828 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1829 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1830 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1831 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1832 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1833 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1834 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1835 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1836 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1837 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1838 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1839 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1840 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1841 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1842 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1843 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1844 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1845 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1846 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1847 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1848 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1849 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1850 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1851 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1852 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1853 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1854 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1855 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1856 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1857 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1858 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1859 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1860 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1861 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1862 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1863 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1864 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1865 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1866 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1867 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1868 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1869 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1870 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1871 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1872 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1873 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1874 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1875 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1876 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1877 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1878 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1879 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1880 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1881 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1882 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1883 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1884 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1885 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1886 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1887 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1888 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1889 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1890 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1891 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1892 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1893 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1894 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1895 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1896 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1897 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1898 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1899 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1900 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1901 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1902 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		others => x"00000000"
	);


begin

	process(i_clk)
	begin
		if rising_edge(i_clk) then
			-- memory write --
			if i_we = '1' then
				mem(to_integer(unsigned(i_w_addr))) <= i_data;
			end if;
			-- memory read -- 
			o_data <= mem(to_integer(unsigned(i_r_addr)));
			
		end if; 
	end process;

end architecture arch;